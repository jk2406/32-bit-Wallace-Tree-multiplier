VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wallacetree32x32
  CLASS BLOCK ;
  FOREIGN wallacetree32x32 ;
  ORIGIN 0.000 0.000 ;
  SIZE 416.055 BY 426.775 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 413.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 413.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.540 10.640 333.140 413.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 30.030 410.560 31.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 183.210 410.560 184.810 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 336.390 410.560 337.990 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 413.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 413.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 413.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.730 410.560 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 179.910 410.560 181.510 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 333.090 410.560 334.690 ;
    END
  END VPWR
  PIN a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 412.055 414.840 416.055 415.440 ;
    END
  END a[0]
  PIN a[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 412.055 156.440 416.055 157.040 ;
    END
  END a[10]
  PIN a[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 412.055 238.040 416.055 238.640 ;
    END
  END a[11]
  PIN a[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 336.640 4.000 337.240 ;
    END
  END a[12]
  PIN a[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 183.630 422.775 183.910 426.775 ;
    END
  END a[13]
  PIN a[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.040 4.000 323.640 ;
    END
  END a[14]
  PIN a[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 196.510 422.775 196.790 426.775 ;
    END
  END a[15]
  PIN a[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 296.330 0.000 296.610 4.000 ;
    END
  END a[16]
  PIN a[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END a[17]
  PIN a[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 351.070 422.775 351.350 426.775 ;
    END
  END a[18]
  PIN a[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 67.710 422.775 67.990 426.775 ;
    END
  END a[19]
  PIN a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 363.950 422.775 364.230 426.775 ;
    END
  END a[1]
  PIN a[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 412.250 0.000 412.530 4.000 ;
    END
  END a[20]
  PIN a[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END a[21]
  PIN a[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END a[22]
  PIN a[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 412.055 142.840 416.055 143.440 ;
    END
  END a[23]
  PIN a[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 415.470 422.775 415.750 426.775 ;
    END
  END a[24]
  PIN a[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 412.055 102.040 416.055 102.640 ;
    END
  END a[25]
  PIN a[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END a[26]
  PIN a[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 170.750 422.775 171.030 426.775 ;
    END
  END a[27]
  PIN a[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 412.055 319.640 416.055 320.240 ;
    END
  END a[28]
  PIN a[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END a[29]
  PIN a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END a[2]
  PIN a[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 93.470 422.775 93.750 426.775 ;
    END
  END a[30]
  PIN a[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 412.055 251.640 416.055 252.240 ;
    END
  END a[31]
  PIN a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END a[3]
  PIN a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 389.710 422.775 389.990 426.775 ;
    END
  END a[4]
  PIN a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 222.270 422.775 222.550 426.775 ;
    END
  END a[5]
  PIN a[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 412.055 292.440 416.055 293.040 ;
    END
  END a[6]
  PIN a[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 260.910 422.775 261.190 426.775 ;
    END
  END a[7]
  PIN a[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 399.370 0.000 399.650 4.000 ;
    END
  END a[8]
  PIN a[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 412.055 210.840 416.055 211.440 ;
    END
  END a[9]
  PIN b[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.840 4.000 296.440 ;
    END
  END b[0]
  PIN b[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 412.055 306.040 416.055 306.640 ;
    END
  END b[10]
  PIN b[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END b[11]
  PIN b[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 402.590 422.775 402.870 426.775 ;
    END
  END b[12]
  PIN b[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 347.850 0.000 348.130 4.000 ;
    END
  END b[13]
  PIN b[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 322.090 0.000 322.370 4.000 ;
    END
  END b[14]
  PIN b[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END b[15]
  PIN b[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END b[16]
  PIN b[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END b[17]
  PIN b[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END b[18]
  PIN b[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 235.150 422.775 235.430 426.775 ;
    END
  END b[19]
  PIN b[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END b[1]
  PIN b[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.240 4.000 214.840 ;
    END
  END b[20]
  PIN b[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 41.950 422.775 42.230 426.775 ;
    END
  END b[21]
  PIN b[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 286.670 422.775 286.950 426.775 ;
    END
  END b[22]
  PIN b[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 119.230 422.775 119.510 426.775 ;
    END
  END b[23]
  PIN b[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.040 4.000 255.640 ;
    END
  END b[24]
  PIN b[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END b[25]
  PIN b[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END b[26]
  PIN b[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 412.055 34.040 416.055 34.640 ;
    END
  END b[27]
  PIN b[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 4.000 ;
    END
  END b[28]
  PIN b[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END b[29]
  PIN b[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 412.055 401.240 416.055 401.840 ;
    END
  END b[2]
  PIN b[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.240 4.000 418.840 ;
    END
  END b[30]
  PIN b[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END b[31]
  PIN b[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 106.350 422.775 106.630 426.775 ;
    END
  END b[3]
  PIN b[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.640 4.000 269.240 ;
    END
  END b[4]
  PIN b[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 412.055 374.040 416.055 374.640 ;
    END
  END b[5]
  PIN b[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 412.055 333.240 416.055 333.840 ;
    END
  END b[6]
  PIN b[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 29.070 422.775 29.350 426.775 ;
    END
  END b[7]
  PIN b[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 54.830 422.775 55.110 426.775 ;
    END
  END b[8]
  PIN b[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END b[9]
  PIN prod[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END prod[0]
  PIN prod[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 144.990 422.775 145.270 426.775 ;
    END
  END prod[10]
  PIN prod[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 412.055 170.040 416.055 170.640 ;
    END
  END prod[11]
  PIN prod[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 412.055 115.640 416.055 116.240 ;
    END
  END prod[12]
  PIN prod[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 309.440 4.000 310.040 ;
    END
  END prod[13]
  PIN prod[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 157.870 422.775 158.150 426.775 ;
    END
  END prod[14]
  PIN prod[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 412.055 6.840 416.055 7.440 ;
    END
  END prod[15]
  PIN prod[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 412.055 129.240 416.055 129.840 ;
    END
  END prod[16]
  PIN prod[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 325.310 422.775 325.590 426.775 ;
    END
  END prod[17]
  PIN prod[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 412.055 74.840 416.055 75.440 ;
    END
  END prod[18]
  PIN prod[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 360.730 0.000 361.010 4.000 ;
    END
  END prod[19]
  PIN prod[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 241.440 4.000 242.040 ;
    END
  END prod[1]
  PIN prod[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END prod[20]
  PIN prod[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 412.055 387.640 416.055 388.240 ;
    END
  END prod[21]
  PIN prod[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END prod[22]
  PIN prod[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 412.055 47.640 416.055 48.240 ;
    END
  END prod[23]
  PIN prod[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.040 4.000 391.640 ;
    END
  END prod[24]
  PIN prod[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 386.490 0.000 386.770 4.000 ;
    END
  END prod[25]
  PIN prod[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 209.390 422.775 209.670 426.775 ;
    END
  END prod[26]
  PIN prod[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END prod[27]
  PIN prod[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END prod[28]
  PIN prod[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END prod[29]
  PIN prod[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 412.055 20.440 416.055 21.040 ;
    END
  END prod[2]
  PIN prod[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END prod[30]
  PIN prod[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 412.055 183.640 416.055 184.240 ;
    END
  END prod[31]
  PIN prod[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 334.970 0.000 335.250 4.000 ;
    END
  END prod[32]
  PIN prod[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.240 4.000 282.840 ;
    END
  END prod[33]
  PIN prod[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 412.055 88.440 416.055 89.040 ;
    END
  END prod[34]
  PIN prod[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 377.440 4.000 378.040 ;
    END
  END prod[35]
  PIN prod[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 412.055 224.440 416.055 225.040 ;
    END
  END prod[36]
  PIN prod[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 412.055 346.840 416.055 347.440 ;
    END
  END prod[37]
  PIN prod[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 373.610 0.000 373.890 4.000 ;
    END
  END prod[38]
  PIN prod[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 412.055 360.440 416.055 361.040 ;
    END
  END prod[39]
  PIN prod[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END prod[3]
  PIN prod[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 4.000 201.240 ;
    END
  END prod[40]
  PIN prod[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END prod[41]
  PIN prod[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END prod[42]
  PIN prod[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 270.570 0.000 270.850 4.000 ;
    END
  END prod[43]
  PIN prod[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 3.310 422.775 3.590 426.775 ;
    END
  END prod[44]
  PIN prod[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 132.110 422.775 132.390 426.775 ;
    END
  END prod[45]
  PIN prod[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 273.790 422.775 274.070 426.775 ;
    END
  END prod[46]
  PIN prod[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.240 4.000 350.840 ;
    END
  END prod[47]
  PIN prod[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.440 4.000 174.040 ;
    END
  END prod[48]
  PIN prod[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END prod[49]
  PIN prod[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 338.190 422.775 338.470 426.775 ;
    END
  END prod[4]
  PIN prod[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 248.030 422.775 248.310 426.775 ;
    END
  END prod[50]
  PIN prod[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END prod[51]
  PIN prod[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 376.830 422.775 377.110 426.775 ;
    END
  END prod[52]
  PIN prod[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 412.055 61.240 416.055 61.840 ;
    END
  END prod[53]
  PIN prod[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 404.640 4.000 405.240 ;
    END
  END prod[54]
  PIN prod[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 412.055 265.240 416.055 265.840 ;
    END
  END prod[55]
  PIN prod[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END prod[56]
  PIN prod[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END prod[57]
  PIN prod[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END prod[58]
  PIN prod[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 412.055 278.840 416.055 279.440 ;
    END
  END prod[59]
  PIN prod[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 4.000 ;
    END
  END prod[5]
  PIN prod[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 312.430 422.775 312.710 426.775 ;
    END
  END prod[60]
  PIN prod[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 299.550 422.775 299.830 426.775 ;
    END
  END prod[61]
  PIN prod[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 16.190 422.775 16.470 426.775 ;
    END
  END prod[62]
  PIN prod[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 80.590 422.775 80.870 426.775 ;
    END
  END prod[63]
  PIN prod[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 283.450 0.000 283.730 4.000 ;
    END
  END prod[6]
  PIN prod[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END prod[7]
  PIN prod[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.840 4.000 364.440 ;
    END
  END prod[8]
  PIN prod[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 412.055 197.240 416.055 197.840 ;
    END
  END prod[9]
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 410.320 413.525 ;
      LAYER met1 ;
        RECT 0.070 9.560 415.770 413.680 ;
      LAYER met2 ;
        RECT 0.100 422.495 3.030 423.370 ;
        RECT 3.870 422.495 15.910 423.370 ;
        RECT 16.750 422.495 28.790 423.370 ;
        RECT 29.630 422.495 41.670 423.370 ;
        RECT 42.510 422.495 54.550 423.370 ;
        RECT 55.390 422.495 67.430 423.370 ;
        RECT 68.270 422.495 80.310 423.370 ;
        RECT 81.150 422.495 93.190 423.370 ;
        RECT 94.030 422.495 106.070 423.370 ;
        RECT 106.910 422.495 118.950 423.370 ;
        RECT 119.790 422.495 131.830 423.370 ;
        RECT 132.670 422.495 144.710 423.370 ;
        RECT 145.550 422.495 157.590 423.370 ;
        RECT 158.430 422.495 170.470 423.370 ;
        RECT 171.310 422.495 183.350 423.370 ;
        RECT 184.190 422.495 196.230 423.370 ;
        RECT 197.070 422.495 209.110 423.370 ;
        RECT 209.950 422.495 221.990 423.370 ;
        RECT 222.830 422.495 234.870 423.370 ;
        RECT 235.710 422.495 247.750 423.370 ;
        RECT 248.590 422.495 260.630 423.370 ;
        RECT 261.470 422.495 273.510 423.370 ;
        RECT 274.350 422.495 286.390 423.370 ;
        RECT 287.230 422.495 299.270 423.370 ;
        RECT 300.110 422.495 312.150 423.370 ;
        RECT 312.990 422.495 325.030 423.370 ;
        RECT 325.870 422.495 337.910 423.370 ;
        RECT 338.750 422.495 350.790 423.370 ;
        RECT 351.630 422.495 363.670 423.370 ;
        RECT 364.510 422.495 376.550 423.370 ;
        RECT 377.390 422.495 389.430 423.370 ;
        RECT 390.270 422.495 402.310 423.370 ;
        RECT 403.150 422.495 415.190 423.370 ;
        RECT 0.100 4.280 415.740 422.495 ;
        RECT 0.650 4.000 12.690 4.280 ;
        RECT 13.530 4.000 25.570 4.280 ;
        RECT 26.410 4.000 38.450 4.280 ;
        RECT 39.290 4.000 51.330 4.280 ;
        RECT 52.170 4.000 64.210 4.280 ;
        RECT 65.050 4.000 77.090 4.280 ;
        RECT 77.930 4.000 89.970 4.280 ;
        RECT 90.810 4.000 102.850 4.280 ;
        RECT 103.690 4.000 115.730 4.280 ;
        RECT 116.570 4.000 128.610 4.280 ;
        RECT 129.450 4.000 141.490 4.280 ;
        RECT 142.330 4.000 154.370 4.280 ;
        RECT 155.210 4.000 167.250 4.280 ;
        RECT 168.090 4.000 180.130 4.280 ;
        RECT 180.970 4.000 193.010 4.280 ;
        RECT 193.850 4.000 205.890 4.280 ;
        RECT 206.730 4.000 218.770 4.280 ;
        RECT 219.610 4.000 231.650 4.280 ;
        RECT 232.490 4.000 244.530 4.280 ;
        RECT 245.370 4.000 257.410 4.280 ;
        RECT 258.250 4.000 270.290 4.280 ;
        RECT 271.130 4.000 283.170 4.280 ;
        RECT 284.010 4.000 296.050 4.280 ;
        RECT 296.890 4.000 308.930 4.280 ;
        RECT 309.770 4.000 321.810 4.280 ;
        RECT 322.650 4.000 334.690 4.280 ;
        RECT 335.530 4.000 347.570 4.280 ;
        RECT 348.410 4.000 360.450 4.280 ;
        RECT 361.290 4.000 373.330 4.280 ;
        RECT 374.170 4.000 386.210 4.280 ;
        RECT 387.050 4.000 399.090 4.280 ;
        RECT 399.930 4.000 411.970 4.280 ;
        RECT 412.810 4.000 415.740 4.280 ;
      LAYER met3 ;
        RECT 4.400 417.840 412.055 418.705 ;
        RECT 3.990 415.840 412.055 417.840 ;
        RECT 3.990 414.440 411.655 415.840 ;
        RECT 3.990 405.640 412.055 414.440 ;
        RECT 4.400 404.240 412.055 405.640 ;
        RECT 3.990 402.240 412.055 404.240 ;
        RECT 3.990 400.840 411.655 402.240 ;
        RECT 3.990 392.040 412.055 400.840 ;
        RECT 4.400 390.640 412.055 392.040 ;
        RECT 3.990 388.640 412.055 390.640 ;
        RECT 3.990 387.240 411.655 388.640 ;
        RECT 3.990 378.440 412.055 387.240 ;
        RECT 4.400 377.040 412.055 378.440 ;
        RECT 3.990 375.040 412.055 377.040 ;
        RECT 3.990 373.640 411.655 375.040 ;
        RECT 3.990 364.840 412.055 373.640 ;
        RECT 4.400 363.440 412.055 364.840 ;
        RECT 3.990 361.440 412.055 363.440 ;
        RECT 3.990 360.040 411.655 361.440 ;
        RECT 3.990 351.240 412.055 360.040 ;
        RECT 4.400 349.840 412.055 351.240 ;
        RECT 3.990 347.840 412.055 349.840 ;
        RECT 3.990 346.440 411.655 347.840 ;
        RECT 3.990 337.640 412.055 346.440 ;
        RECT 4.400 336.240 412.055 337.640 ;
        RECT 3.990 334.240 412.055 336.240 ;
        RECT 3.990 332.840 411.655 334.240 ;
        RECT 3.990 324.040 412.055 332.840 ;
        RECT 4.400 322.640 412.055 324.040 ;
        RECT 3.990 320.640 412.055 322.640 ;
        RECT 3.990 319.240 411.655 320.640 ;
        RECT 3.990 310.440 412.055 319.240 ;
        RECT 4.400 309.040 412.055 310.440 ;
        RECT 3.990 307.040 412.055 309.040 ;
        RECT 3.990 305.640 411.655 307.040 ;
        RECT 3.990 296.840 412.055 305.640 ;
        RECT 4.400 295.440 412.055 296.840 ;
        RECT 3.990 293.440 412.055 295.440 ;
        RECT 3.990 292.040 411.655 293.440 ;
        RECT 3.990 283.240 412.055 292.040 ;
        RECT 4.400 281.840 412.055 283.240 ;
        RECT 3.990 279.840 412.055 281.840 ;
        RECT 3.990 278.440 411.655 279.840 ;
        RECT 3.990 269.640 412.055 278.440 ;
        RECT 4.400 268.240 412.055 269.640 ;
        RECT 3.990 266.240 412.055 268.240 ;
        RECT 3.990 264.840 411.655 266.240 ;
        RECT 3.990 256.040 412.055 264.840 ;
        RECT 4.400 254.640 412.055 256.040 ;
        RECT 3.990 252.640 412.055 254.640 ;
        RECT 3.990 251.240 411.655 252.640 ;
        RECT 3.990 242.440 412.055 251.240 ;
        RECT 4.400 241.040 412.055 242.440 ;
        RECT 3.990 239.040 412.055 241.040 ;
        RECT 3.990 237.640 411.655 239.040 ;
        RECT 3.990 228.840 412.055 237.640 ;
        RECT 4.400 227.440 412.055 228.840 ;
        RECT 3.990 225.440 412.055 227.440 ;
        RECT 3.990 224.040 411.655 225.440 ;
        RECT 3.990 215.240 412.055 224.040 ;
        RECT 4.400 213.840 412.055 215.240 ;
        RECT 3.990 211.840 412.055 213.840 ;
        RECT 3.990 210.440 411.655 211.840 ;
        RECT 3.990 201.640 412.055 210.440 ;
        RECT 4.400 200.240 412.055 201.640 ;
        RECT 3.990 198.240 412.055 200.240 ;
        RECT 3.990 196.840 411.655 198.240 ;
        RECT 3.990 188.040 412.055 196.840 ;
        RECT 4.400 186.640 412.055 188.040 ;
        RECT 3.990 184.640 412.055 186.640 ;
        RECT 3.990 183.240 411.655 184.640 ;
        RECT 3.990 174.440 412.055 183.240 ;
        RECT 4.400 173.040 412.055 174.440 ;
        RECT 3.990 171.040 412.055 173.040 ;
        RECT 3.990 169.640 411.655 171.040 ;
        RECT 3.990 160.840 412.055 169.640 ;
        RECT 4.400 159.440 412.055 160.840 ;
        RECT 3.990 157.440 412.055 159.440 ;
        RECT 3.990 156.040 411.655 157.440 ;
        RECT 3.990 147.240 412.055 156.040 ;
        RECT 4.400 145.840 412.055 147.240 ;
        RECT 3.990 143.840 412.055 145.840 ;
        RECT 3.990 142.440 411.655 143.840 ;
        RECT 3.990 133.640 412.055 142.440 ;
        RECT 4.400 132.240 412.055 133.640 ;
        RECT 3.990 130.240 412.055 132.240 ;
        RECT 3.990 128.840 411.655 130.240 ;
        RECT 3.990 120.040 412.055 128.840 ;
        RECT 4.400 118.640 412.055 120.040 ;
        RECT 3.990 116.640 412.055 118.640 ;
        RECT 3.990 115.240 411.655 116.640 ;
        RECT 3.990 106.440 412.055 115.240 ;
        RECT 4.400 105.040 412.055 106.440 ;
        RECT 3.990 103.040 412.055 105.040 ;
        RECT 3.990 101.640 411.655 103.040 ;
        RECT 3.990 92.840 412.055 101.640 ;
        RECT 4.400 91.440 412.055 92.840 ;
        RECT 3.990 89.440 412.055 91.440 ;
        RECT 3.990 88.040 411.655 89.440 ;
        RECT 3.990 79.240 412.055 88.040 ;
        RECT 4.400 77.840 412.055 79.240 ;
        RECT 3.990 75.840 412.055 77.840 ;
        RECT 3.990 74.440 411.655 75.840 ;
        RECT 3.990 65.640 412.055 74.440 ;
        RECT 4.400 64.240 412.055 65.640 ;
        RECT 3.990 62.240 412.055 64.240 ;
        RECT 3.990 60.840 411.655 62.240 ;
        RECT 3.990 52.040 412.055 60.840 ;
        RECT 4.400 50.640 412.055 52.040 ;
        RECT 3.990 48.640 412.055 50.640 ;
        RECT 3.990 47.240 411.655 48.640 ;
        RECT 3.990 38.440 412.055 47.240 ;
        RECT 4.400 37.040 412.055 38.440 ;
        RECT 3.990 35.040 412.055 37.040 ;
        RECT 3.990 33.640 411.655 35.040 ;
        RECT 3.990 24.840 412.055 33.640 ;
        RECT 4.400 23.440 412.055 24.840 ;
        RECT 3.990 21.440 412.055 23.440 ;
        RECT 3.990 20.040 411.655 21.440 ;
        RECT 3.990 11.240 412.055 20.040 ;
        RECT 4.400 9.840 412.055 11.240 ;
        RECT 3.990 7.840 412.055 9.840 ;
        RECT 3.990 6.975 411.655 7.840 ;
      LAYER met4 ;
        RECT 40.775 13.095 174.240 411.905 ;
        RECT 176.640 13.095 177.540 411.905 ;
        RECT 179.940 13.095 327.840 411.905 ;
        RECT 330.240 13.095 331.140 411.905 ;
        RECT 333.540 13.095 381.505 411.905 ;
      LAYER met5 ;
        RECT 279.340 164.100 344.420 165.700 ;
  END
END wallacetree32x32
END LIBRARY

