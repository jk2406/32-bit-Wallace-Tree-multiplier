* NGSPICE file created from wallacetree32x32.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_4 abstract view
.subckt sky130_fd_sc_hd__o2111a_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_4 abstract view
.subckt sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd1_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd1_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_4 abstract view
.subckt sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_4 abstract view
.subckt sky130_fd_sc_hd__o21ba_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_4 abstract view
.subckt sky130_fd_sc_hd__nor2b_4 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_2 abstract view
.subckt sky130_fd_sc_hd__o32ai_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_4 abstract view
.subckt sky130_fd_sc_hd__o41a_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_4 abstract view
.subckt sky130_fd_sc_hd__a41oi_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_4 abstract view
.subckt sky130_fd_sc_hd__or2b_4 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_4 abstract view
.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s4s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s4s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_4 abstract view
.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_4 abstract view
.subckt sky130_fd_sc_hd__a2111oi_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

.subckt wallacetree32x32 VGND VPWR a[0] a[10] a[11] a[12] a[13] a[14] a[15] a[16]
+ a[17] a[18] a[19] a[1] a[20] a[21] a[22] a[23] a[24] a[25] a[26] a[27] a[28] a[29]
+ a[2] a[30] a[31] a[3] a[4] a[5] a[6] a[7] a[8] a[9] b[0] b[10] b[11] b[12] b[13]
+ b[14] b[15] b[16] b[17] b[18] b[19] b[1] b[20] b[21] b[22] b[23] b[24] b[25] b[26]
+ b[27] b[28] b[29] b[2] b[30] b[31] b[3] b[4] b[5] b[6] b[7] b[8] b[9] prod[0] prod[10]
+ prod[11] prod[12] prod[13] prod[14] prod[15] prod[16] prod[17] prod[18] prod[19]
+ prod[1] prod[20] prod[21] prod[22] prod[23] prod[24] prod[25] prod[26] prod[27]
+ prod[28] prod[29] prod[2] prod[30] prod[31] prod[32] prod[33] prod[34] prod[35]
+ prod[36] prod[37] prod[38] prod[39] prod[3] prod[40] prod[41] prod[42] prod[43]
+ prod[44] prod[45] prod[46] prod[47] prod[48] prod[49] prod[4] prod[50] prod[51]
+ prod[52] prod[53] prod[54] prod[55] prod[56] prod[57] prod[58] prod[59] prod[5]
+ prod[60] prod[61] prod[62] prod[63] prod[6] prod[7] prod[8] prod[9]
XANTENNA__10669__A1 _05181_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09671_ _01724_ _01726_ _01846_ VGND VGND VPWR VPWR _01848_ sky130_fd_sc_hd__nor3_1
X_08622_ _00699_ _00700_ VGND VGND VPWR VPWR _00701_ sky130_fd_sc_hd__nor2_2
X_08553_ _00623_ _00609_ _00610_ VGND VGND VPWR VPWR _00625_ sky130_fd_sc_hd__and3_1
XFILLER_0_76_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07504_ _04862_ VGND VGND VPWR VPWR _04895_ sky130_fd_sc_hd__clkbuf_4
X_08484_ _00465_ _00548_ _00549_ VGND VGND VPWR VPWR _00550_ sky130_fd_sc_hd__nor3_1
XFILLER_0_134_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07435_ _04114_ _04125_ VGND VGND VPWR VPWR _04136_ sky130_fd_sc_hd__and2b_1
XFILLER_0_64_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10974__A _04917_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07366_ _03356_ net188 VGND VGND VPWR VPWR _03378_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_91_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11397__A2 _01254_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09105_ _00530_ _00391_ _01228_ VGND VGND VPWR VPWR _01229_ sky130_fd_sc_hd__and3_1
XFILLER_0_115_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07297_ _02598_ _02609_ VGND VGND VPWR VPWR _02620_ sky130_fd_sc_hd__and2b_1
XANTENNA__13500__D _03680_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09036_ _01117_ _01151_ _01118_ VGND VGND VPWR VPWR _01154_ sky130_fd_sc_hd__nor3_1
XFILLER_0_130_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09275__A _01414_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09938_ _02132_ _02140_ VGND VGND VPWR VPWR _02141_ sky130_fd_sc_hd__xor2_1
X_09869_ _06964_ _00121_ _00755_ _00741_ VGND VGND VPWR VPWR _02065_ sky130_fd_sc_hd__nand4_2
XFILLER_0_99_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11900_ _02040_ _03681_ _04144_ _04143_ _02135_ VGND VGND VPWR VPWR _04295_ sky130_fd_sc_hd__a32o_1
XTAP_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12880_ _00605_ _02120_ VGND VGND VPWR VPWR _05373_ sky130_fd_sc_hd__nand2_1
XTAP_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11609__B1 _01250_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11831_ _02660_ _04218_ VGND VGND VPWR VPWR _04219_ sky130_fd_sc_hd__xnor2_1
XTAP_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09441__C _00574_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07828__A2 net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11762_ _00138_ _02018_ _01953_ VGND VGND VPWR VPWR _04143_ sky130_fd_sc_hd__and3_1
XFILLER_0_138_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13501_ _01415_ _03680_ _06035_ _06036_ VGND VGND VPWR VPWR _06038_ sky130_fd_sc_hd__o2bb2a_1
X_10713_ _02937_ _02939_ _02948_ _02989_ VGND VGND VPWR VPWR _02990_ sky130_fd_sc_hd__or4_1
XFILLER_0_95_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11693_ _04065_ _04066_ VGND VGND VPWR VPWR _04067_ sky130_fd_sc_hd__nor2_1
XTAP_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13432_ _05628_ _05630_ _05421_ VGND VGND VPWR VPWR _05963_ sky130_fd_sc_hd__a21o_1
X_10644_ _02903_ _02912_ VGND VGND VPWR VPWR _02914_ sky130_fd_sc_hd__or2_1
XANTENNA__08354__A _00395_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12585__A1 _03740_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12585__B2 _03707_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10575_ _02835_ _02837_ VGND VGND VPWR VPWR _02838_ sky130_fd_sc_hd__nor2_1
X_13363_ _00416_ _01288_ _02720_ VGND VGND VPWR VPWR _05887_ sky130_fd_sc_hd__and3_1
XFILLER_0_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer7 _00825_ VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__buf_1
XFILLER_0_106_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12314_ _00459_ _01780_ _04749_ VGND VGND VPWR VPWR _04750_ sky130_fd_sc_hd__and3_1
XFILLER_0_133_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_411 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13294_ _05798_ _05815_ VGND VGND VPWR VPWR _05816_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_792 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12245_ _00783_ _01178_ _01248_ _04037_ VGND VGND VPWR VPWR _04674_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12176_ _04018_ _04019_ VGND VGND VPWR VPWR _04599_ sky130_fd_sc_hd__nand2_1
XANTENNA__09653__C_N _01828_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11127_ _03369_ _03384_ _03443_ VGND VGND VPWR VPWR _03446_ sky130_fd_sc_hd__o21a_1
X_11058_ _03365_ _03368_ VGND VGND VPWR VPWR _03370_ sky130_fd_sc_hd__nor2_1
XANTENNA__09913__A _02007_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10009_ _02211_ _02217_ VGND VGND VPWR VPWR _02219_ sky130_fd_sc_hd__nand2_1
XANTENNA__07433__A _03576_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07152__B net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10823__A1 _01339_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07220_ _01656_ _01667_ VGND VGND VPWR VPWR _01777_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_144_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08264__A _02040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_715 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11902__A2_N _03682_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07151_ _00967_ _01011_ VGND VGND VPWR VPWR _01022_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10960__C _02187_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11000__A1 _04378_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11000__B2 _02971_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10034__A _00843_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13828__A1 _04714_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07984_ _00026_ _00027_ VGND VGND VPWR VPWR _00028_ sky130_fd_sc_hd__or2_1
X_09723_ _01890_ _01903_ VGND VGND VPWR VPWR _01905_ sky130_fd_sc_hd__nor2_1
XANTENNA__09823__A _06818_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11839__B1 _03686_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12500__A1 _00612_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12500__B2 _04026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09654_ _01759_ _01760_ _01828_ VGND VGND VPWR VPWR _01830_ sky130_fd_sc_hd__o21bai_2
XANTENNA__11791__C _01744_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10688__B _02982_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08605_ _00678_ _00680_ VGND VGND VPWR VPWR _00682_ sky130_fd_sc_hd__and2_1
XANTENNA__13056__A2 _02703_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09585_ _01443_ _01444_ _01753_ VGND VGND VPWR VPWR _01754_ sky130_fd_sc_hd__a21o_1
XFILLER_0_145_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08536_ _00605_ VGND VGND VPWR VPWR _00607_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08467_ _02993_ _06873_ _06875_ _05203_ VGND VGND VPWR VPWR _00532_ sky130_fd_sc_hd__and4_1
XFILLER_0_65_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07418_ _00311_ _03938_ VGND VGND VPWR VPWR _03949_ sky130_fd_sc_hd__nand2_1
X_08398_ _00454_ _00455_ VGND VGND VPWR VPWR _00456_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_512 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07349_ _03136_ _03180_ VGND VGND VPWR VPWR _03191_ sky130_fd_sc_hd__xor2_1
XFILLER_0_73_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10360_ _06733_ _03773_ VGND VGND VPWR VPWR _02603_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_578 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09019_ _06965_ _04906_ VGND VGND VPWR VPWR _01135_ sky130_fd_sc_hd__nand2_1
XANTENNA__11790__A2 _02133_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10291_ _05577_ _01410_ VGND VGND VPWR VPWR _02527_ sky130_fd_sc_hd__nand2_1
XFILLER_0_131_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12030_ _04436_ _04437_ VGND VGND VPWR VPWR _04438_ sky130_fd_sc_hd__nor2_1
XFILLER_0_103_488 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13819__A1 _02187_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13819__B2 _01400_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13981_ _06550_ _06552_ VGND VGND VPWR VPWR _06566_ sky130_fd_sc_hd__and2_1
XANTENNA__13255__A _05524_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12932_ _05426_ _05429_ VGND VGND VPWR VPWR _05430_ sky130_fd_sc_hd__xor2_2
XFILLER_0_88_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07253__A _02127_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12863_ _05275_ _05293_ VGND VGND VPWR VPWR _05354_ sky130_fd_sc_hd__nand2_1
XTAP_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13405__D _03686_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11814_ _04198_ _04194_ _04195_ VGND VGND VPWR VPWR _04200_ sky130_fd_sc_hd__nor3_1
XTAP_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12794_ _00914_ _02168_ VGND VGND VPWR VPWR _05278_ sky130_fd_sc_hd__nand2_1
XTAP_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11745_ _04119_ _04123_ VGND VGND VPWR VPWR _04124_ sky130_fd_sc_hd__xor2_1
XTAP_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11676_ _00112_ _00268_ _00755_ _01260_ VGND VGND VPWR VPWR _04049_ sky130_fd_sc_hd__nand4_1
XFILLER_0_24_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_512 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13415_ _05898_ _05942_ VGND VGND VPWR VPWR _05944_ sky130_fd_sc_hd__or2_1
X_10627_ _02805_ _02812_ VGND VGND VPWR VPWR _02896_ sky130_fd_sc_hd__and2b_1
XANTENNA__08226__A2 _00112_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_843 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09423__A1 _06417_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13346_ _05340_ _05348_ VGND VGND VPWR VPWR _05869_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10558_ _00293_ _02169_ VGND VGND VPWR VPWR _02820_ sky130_fd_sc_hd__nand2_1
XFILLER_0_106_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13277_ _05604_ _05732_ VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__xnor2_1
XFILLER_0_121_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10489_ _01473_ _02743_ VGND VGND VPWR VPWR _02744_ sky130_fd_sc_hd__nand2_1
XANTENNA__07428__A _04048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12228_ _04652_ _04654_ _04655_ VGND VGND VPWR VPWR _04656_ sky130_fd_sc_hd__and3_1
XANTENNA__07737__A1 _00420_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07737__B2 net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12159_ _02476_ _02480_ _04577_ _04578_ _04579_ VGND VGND VPWR VPWR _04580_ sky130_fd_sc_hd__o2111a_4
XANTENNA__10789__A _00628_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09362__B _01505_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08259__A _06417_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13501__A1_N _01415_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09370_ _06461_ _01518_ VGND VGND VPWR VPWR _01519_ sky130_fd_sc_hd__nand2_1
XANTENNA__12797__A1 _00914_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08321_ _00350_ _00371_ VGND VGND VPWR VPWR _00372_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08252_ _00050_ _00153_ _00292_ _00295_ VGND VGND VPWR VPWR _00296_ sky130_fd_sc_hd__a211o_1
XFILLER_0_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07203_ _00420_ _01208_ _00661_ _00978_ VGND VGND VPWR VPWR _01591_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08183_ _00217_ _00219_ VGND VGND VPWR VPWR _00227_ sky130_fd_sc_hd__xor2_1
XFILLER_0_132_506 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_331 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07134_ _00694_ _00814_ VGND VGND VPWR VPWR _00836_ sky130_fd_sc_hd__nand2_1
XANTENNA__09818__A _00486_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09965__A2 _01934_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10971__B _00457_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09537__B _04026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07338__A _03059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07967_ _00891_ _01120_ _07010_ net38 VGND VGND VPWR VPWR _00011_ sky130_fd_sc_hd__nand4_1
X_09706_ _01883_ _01884_ VGND VGND VPWR VPWR _01887_ sky130_fd_sc_hd__or2_1
X_07898_ _07021_ _07026_ VGND VGND VPWR VPWR _07027_ sky130_fd_sc_hd__xor2_1
XANTENNA__08906__A2_N _00095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10849__D net52 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09637_ _01744_ net19 VGND VGND VPWR VPWR _01812_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13803__A _03414_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09568_ _01476_ _01734_ VGND VGND VPWR VPWR _01736_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08519_ _03982_ _00430_ _00429_ VGND VGND VPWR VPWR _00588_ sky130_fd_sc_hd__a21boi_2
X_09499_ _01654_ _01659_ VGND VGND VPWR VPWR _01660_ sky130_fd_sc_hd__xor2_1
XFILLER_0_77_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11530_ _03884_ _03886_ _03887_ VGND VGND VPWR VPWR _03888_ sky130_fd_sc_hd__a21bo_2
XANTENNA__08781__B1_N _00666_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11042__B _04059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11461_ _03532_ _00121_ _01953_ _02134_ VGND VGND VPWR VPWR _03812_ sky130_fd_sc_hd__nand4_1
XFILLER_0_135_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13200_ _05715_ _05724_ VGND VGND VPWR VPWR _05725_ sky130_fd_sc_hd__xor2_2
XFILLER_0_104_720 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10412_ _02454_ _02659_ VGND VGND VPWR VPWR _02660_ sky130_fd_sc_hd__nor2_1
XFILLER_0_116_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14180_ _02743_ _04014_ _02742_ _04013_ VGND VGND VPWR VPWR _06780_ sky130_fd_sc_hd__and4_1
X_11392_ _00112_ _00268_ _01179_ _01254_ VGND VGND VPWR VPWR _03736_ sky130_fd_sc_hd__and4_1
XFILLER_0_33_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_375 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13131_ _03626_ _03671_ VGND VGND VPWR VPWR _05649_ sky130_fd_sc_hd__xnor2_2
XANTENNA__11763__A2 _01953_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10343_ _02334_ _02345_ VGND VGND VPWR VPWR _02584_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10274_ _00989_ _02312_ net57 _03576_ VGND VGND VPWR VPWR _02508_ sky130_fd_sc_hd__a22o_1
X_13062_ _05568_ _05570_ _05572_ VGND VGND VPWR VPWR _05573_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_29_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12013_ _04408_ _04418_ VGND VGND VPWR VPWR _04419_ sky130_fd_sc_hd__and2b_1
XANTENNA__12304__D _01601_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10105__C net50 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07195__A2 _01197_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13964_ _06535_ _06546_ VGND VGND VPWR VPWR _06547_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08079__A _05566_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09341__B1 _01486_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12915_ _05409_ _05304_ _05410_ VGND VGND VPWR VPWR _05411_ sky130_fd_sc_hd__and3_1
X_13895_ _05937_ _05940_ VGND VGND VPWR VPWR _06471_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12846_ _05286_ _05333_ VGND VGND VPWR VPWR _05336_ sky130_fd_sc_hd__nand2_1
XTAP_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12777_ _04736_ _04773_ VGND VGND VPWR VPWR _05260_ sky130_fd_sc_hd__and2_1
XTAP_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11728_ _04040_ _04105_ VGND VGND VPWR VPWR _04106_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_83_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11659_ _04007_ _03875_ VGND VGND VPWR VPWR _04030_ sky130_fd_sc_hd__and2b_1
XFILLER_0_36_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11203__B2 _03501_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_515 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13329_ _05631_ _05850_ VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__xor2_1
XFILLER_0_110_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12999__A _05487_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08870_ _00776_ _00786_ VGND VGND VPWR VPWR _00972_ sky130_fd_sc_hd__nand2_1
X_07821_ _06862_ _06948_ VGND VGND VPWR VPWR _06950_ sky130_fd_sc_hd__and2_1
XANTENNA__13607__B _03785_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07752_ _06872_ _06880_ VGND VGND VPWR VPWR _06881_ sky130_fd_sc_hd__xnor2_1
X_07683_ net12 net23 net35 net34 VGND VGND VPWR VPWR _06812_ sky130_fd_sc_hd__and4_1
X_09422_ _06428_ _00745_ _01575_ _01263_ VGND VGND VPWR VPWR _01576_ sky130_fd_sc_hd__nand4_1
XFILLER_0_35_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08262__A2_N _00144_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11690__A1 _06819_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11690__B2 _06874_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09353_ _01498_ _01499_ VGND VGND VPWR VPWR _01500_ sky130_fd_sc_hd__or2_2
XFILLER_0_19_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09635__A1 _01197_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09635__B2 _04510_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08436__B _00142_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08304_ _04070_ _04147_ VGND VGND VPWR VPWR _00353_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07340__B _02029_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11442__A1 _06964_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09284_ _01423_ _01424_ VGND VGND VPWR VPWR _01425_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11442__B2 _00121_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_142_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08235_ _00277_ _00278_ VGND VGND VPWR VPWR _00279_ sky130_fd_sc_hd__or2_1
XFILLER_0_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08166_ _06847_ _00209_ VGND VGND VPWR VPWR _00210_ sky130_fd_sc_hd__or2_2
XFILLER_0_43_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07117_ _00639_ VGND VGND VPWR VPWR _00650_ sky130_fd_sc_hd__clkbuf_4
X_08097_ _04917_ _00139_ _00140_ VGND VGND VPWR VPWR _00141_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_113_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13498__A2 _03690_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07218__D _00311_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08999_ _01034_ _01040_ VGND VGND VPWR VPWR _01113_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10579__D _02305_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10961_ _00859_ _02188_ _02190_ _01472_ VGND VGND VPWR VPWR _03263_ sky130_fd_sc_hd__a22oi_1
X_12700_ _05076_ _05077_ VGND VGND VPWR VPWR _05175_ sky130_fd_sc_hd__or2_1
X_13680_ _06201_ _06231_ _06234_ VGND VGND VPWR VPWR _06235_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08627__A _00666_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10892_ _03174_ _03186_ VGND VGND VPWR VPWR _03187_ sky130_fd_sc_hd__nor2_1
XANTENNA__09776__A1_N _01178_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07531__A _04378_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12631_ _05097_ _05098_ VGND VGND VPWR VPWR _05099_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12562_ _00380_ _02008_ _05022_ VGND VGND VPWR VPWR _05023_ sky130_fd_sc_hd__a21o_1
XFILLER_0_53_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11513_ _03715_ _03716_ VGND VGND VPWR VPWR _03869_ sky130_fd_sc_hd__xnor2_4
X_12493_ _00374_ _00755_ _04945_ _04946_ VGND VGND VPWR VPWR _04947_ sky130_fd_sc_hd__a31o_1
XFILLER_0_135_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14232_ _00409_ _00400_ VGND VGND VPWR VPWR _06811_ sky130_fd_sc_hd__or2b_1
X_11444_ _03554_ _03678_ _03791_ _03792_ VGND VGND VPWR VPWR _03793_ sky130_fd_sc_hd__a31o_1
XFILLER_0_22_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08362__A _00415_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14163_ _02742_ _04013_ _06702_ VGND VGND VPWR VPWR _06762_ sky130_fd_sc_hd__and3_1
XFILLER_0_21_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11375_ _03715_ _03716_ VGND VGND VPWR VPWR _03717_ sky130_fd_sc_hd__and2b_1
XFILLER_0_33_194 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13114_ _05315_ _05629_ VGND VGND VPWR VPWR _05630_ sky130_fd_sc_hd__xnor2_2
X_10326_ _04851_ _00780_ _00777_ net4 VGND VGND VPWR VPWR _02566_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14094_ _05821_ _05842_ _06686_ _06687_ _06688_ VGND VGND VPWR VPWR _06689_ sky130_fd_sc_hd__o311a_4
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13045_ _04579_ _05553_ _02701_ VGND VGND VPWR VPWR _05554_ sky130_fd_sc_hd__mux2_4
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13708__A _02427_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10257_ _02279_ _02490_ VGND VGND VPWR VPWR _02491_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_56_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07706__A _00880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10188_ _00486_ _00734_ _02413_ _02414_ VGND VGND VPWR VPWR _02415_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_88_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13947_ _06514_ _06528_ VGND VGND VPWR VPWR _06529_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09640__B net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13878_ _06451_ _06452_ VGND VGND VPWR VPWR _06453_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08537__A _00607_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07441__A _00431_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_423 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12829_ _03675_ VGND VGND VPWR VPWR _05317_ sky130_fd_sc_hd__inv_2
XANTENNA__13162__B _05670_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_724 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_651 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08020_ _00058_ _00063_ VGND VGND VPWR VPWR _00064_ sky130_fd_sc_hd__nor2_1
XFILLER_0_112_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09368__A _00779_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_142_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09971_ _02105_ _02149_ _01058_ _01411_ VGND VGND VPWR VPWR _02177_ sky130_fd_sc_hd__and4_1
XFILLER_0_12_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09560__A2_N _01472_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08922_ _01027_ _01028_ VGND VGND VPWR VPWR _01029_ sky130_fd_sc_hd__or2_1
XANTENNA__07159__A2 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08853_ _00949_ _00952_ VGND VGND VPWR VPWR _00953_ sky130_fd_sc_hd__xor2_1
XFILLER_0_34_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07804_ _04983_ _05291_ VGND VGND VPWR VPWR _06933_ sky130_fd_sc_hd__nand2_1
XANTENNA__07335__B net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08784_ _00553_ _00710_ VGND VGND VPWR VPWR _00878_ sky130_fd_sc_hd__or2_1
X_07735_ _06862_ _06863_ VGND VGND VPWR VPWR _06864_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10977__A _00143_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11663__A1 _00258_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07666_ _06527_ _06648_ VGND VGND VPWR VPWR _06658_ sky130_fd_sc_hd__xor2_2
XFILLER_0_94_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11663__B2 _06765_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09405_ _01493_ _01556_ VGND VGND VPWR VPWR _01557_ sky130_fd_sc_hd__xor2_1
XFILLER_0_48_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13404__A2 _01956_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07597_ _05857_ _05890_ VGND VGND VPWR VPWR _05901_ sky130_fd_sc_hd__nand2_1
X_09336_ _01316_ _01480_ _01345_ VGND VGND VPWR VPWR _01482_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10218__A2 _01177_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13800__B _03682_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09267_ _01064_ _01105_ _01406_ VGND VGND VPWR VPWR _01407_ sky130_fd_sc_hd__and3_1
XFILLER_0_7_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08218_ _06965_ VGND VGND VPWR VPWR _00262_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_90_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09198_ _01134_ _01141_ VGND VGND VPWR VPWR _01331_ sky130_fd_sc_hd__and2_1
XFILLER_0_105_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12416__B _01586_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08149_ _05357_ _00192_ VGND VGND VPWR VPWR _00193_ sky130_fd_sc_hd__nand2_1
XANTENNA__08595__A1 _06472_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08595__B2 _06483_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11160_ _03471_ _03481_ VGND VGND VPWR VPWR _03482_ sky130_fd_sc_hd__nand2_1
XFILLER_0_113_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10111_ _02177_ _02328_ VGND VGND VPWR VPWR _02330_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11091_ _03328_ _03405_ VGND VGND VPWR VPWR _03406_ sky130_fd_sc_hd__nor2_1
X_10042_ _02253_ _02254_ VGND VGND VPWR VPWR _02255_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09741__A _04268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13801_ _02189_ _03686_ _06367_ VGND VGND VPWR VPWR _06368_ sky130_fd_sc_hd__a21boi_1
X_11993_ _04388_ _04391_ _04390_ VGND VGND VPWR VPWR _04397_ sky130_fd_sc_hd__and3_1
X_13732_ _06287_ _06291_ VGND VGND VPWR VPWR _06292_ sky130_fd_sc_hd__nor2_1
X_10944_ _03101_ _03243_ VGND VGND VPWR VPWR _03244_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13663_ _06212_ _06214_ _06215_ VGND VGND VPWR VPWR _06216_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_38_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10875_ _03138_ _03167_ VGND VGND VPWR VPWR _03168_ sky130_fd_sc_hd__and2_1
XFILLER_0_38_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_754 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12614_ _05078_ _05079_ VGND VGND VPWR VPWR _05080_ sky130_fd_sc_hd__nor2_1
X_13594_ _06135_ _06139_ VGND VGND VPWR VPWR _06140_ sky130_fd_sc_hd__and2b_1
XFILLER_0_53_201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12545_ _04816_ VGND VGND VPWR VPWR _05004_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12476_ _04923_ _04927_ VGND VGND VPWR VPWR _04929_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12326__B _02090_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11868__D _01600_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14215_ _03642_ _00229_ VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__xnor2_4
XFILLER_0_34_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11427_ _00004_ _06885_ _01180_ _01249_ VGND VGND VPWR VPWR _03775_ sky130_fd_sc_hd__and4_1
XFILLER_0_22_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14146_ _06714_ _06742_ VGND VGND VPWR VPWR _06745_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_676 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_output86_A net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09916__A _01564_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11358_ _03680_ VGND VGND VPWR VPWR _03699_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08820__A _00157_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13438__A _03785_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10309_ _02353_ _02354_ VGND VGND VPWR VPWR _02547_ sky130_fd_sc_hd__nand2_1
X_14077_ _06668_ _06670_ VGND VGND VPWR VPWR _06671_ sky130_fd_sc_hd__nor2_1
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11289_ _03622_ _03623_ VGND VGND VPWR VPWR _03624_ sky130_fd_sc_hd__and2_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13028_ _04578_ _05535_ VGND VGND VPWR VPWR _05536_ sky130_fd_sc_hd__xnor2_4
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09073__D net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer17 _00182_ VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_83_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrebuffer28 net173 VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer39 _05423_ VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__dlymetal6s2s_1
X_07520_ _04884_ _05049_ VGND VGND VPWR VPWR _05071_ sky130_fd_sc_hd__nand2_1
XANTENNA__09370__B _01518_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07451_ _04158_ _04301_ VGND VGND VPWR VPWR _04312_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07382_ _03543_ VGND VGND VPWR VPWR _03554_ sky130_fd_sc_hd__buf_4
XFILLER_0_146_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09121_ net18 VGND VGND VPWR VPWR _01246_ sky130_fd_sc_hd__buf_2
XFILLER_0_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09052_ _00711_ _00881_ _00882_ _00877_ _01047_ VGND VGND VPWR VPWR _01171_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_115_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08003_ _07045_ _07050_ VGND VGND VPWR VPWR _00047_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_698 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08730__A _00293_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09954_ _01546_ VGND VGND VPWR VPWR _02158_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_110_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12252__A _00378_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08905_ _01008_ _01009_ _06765_ _00095_ VGND VGND VPWR VPWR _01010_ sky130_fd_sc_hd__and4bb_1
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09885_ _02058_ _02081_ VGND VGND VPWR VPWR _02082_ sky130_fd_sc_hd__nor2_1
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08836_ _00932_ _00933_ VGND VGND VPWR VPWR _00935_ sky130_fd_sc_hd__nand2_2
XANTENNA__10687__A2 net50 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08767_ _06626_ _00859_ _00498_ VGND VGND VPWR VPWR _00860_ sky130_fd_sc_hd__and3_1
XFILLER_0_68_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07718_ _06845_ _06846_ VGND VGND VPWR VPWR _06847_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08698_ _00783_ VGND VGND VPWR VPWR _00784_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__07304__A2 _00639_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07649_ _06461_ VGND VGND VPWR VPWR _06472_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_138_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10660_ _02928_ _02930_ _02931_ VGND VGND VPWR VPWR _02932_ sky130_fd_sc_hd__a21o_1
XFILLER_0_94_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09319_ _01461_ _01462_ VGND VGND VPWR VPWR _01463_ sky130_fd_sc_hd__nor2_2
XFILLER_0_91_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10591_ _02855_ VGND VGND VPWR VPWR _02856_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_8_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12330_ _04753_ _04755_ VGND VGND VPWR VPWR _04768_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10611__A2 _01060_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12261_ _04690_ _04691_ VGND VGND VPWR VPWR _04692_ sky130_fd_sc_hd__and2b_1
X_14000_ _06573_ _06578_ _06581_ _06584_ _06586_ VGND VGND VPWR VPWR _06587_ sky130_fd_sc_hd__o311a_1
X_11212_ _03234_ _03237_ VGND VGND VPWR VPWR _03539_ sky130_fd_sc_hd__xor2_1
XANTENNA__13561__B2 _01958_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12192_ _03534_ _03617_ _04615_ VGND VGND VPWR VPWR _04616_ sky130_fd_sc_hd__o21a_1
XANTENNA__10375__A1 _06819_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10375__B2 _06821_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11143_ _03044_ _03029_ _03042_ VGND VGND VPWR VPWR _03463_ sky130_fd_sc_hd__nor3_1
Xoutput75 net75 VGND VGND VPWR VPWR prod[19] sky130_fd_sc_hd__clkbuf_4
Xoutput86 net86 VGND VGND VPWR VPWR prod[29] sky130_fd_sc_hd__clkbuf_4
Xoutput97 net97 VGND VGND VPWR VPWR prod[39] sky130_fd_sc_hd__buf_2
X_11074_ _03382_ _03381_ VGND VGND VPWR VPWR _03387_ sky130_fd_sc_hd__and2b_1
XFILLER_0_37_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10025_ _02209_ _02235_ VGND VGND VPWR VPWR _02236_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_144_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11976_ _04305_ _04314_ _04313_ VGND VGND VPWR VPWR _04379_ sky130_fd_sc_hd__a21oi_1
X_13715_ _02426_ _02759_ _06271_ VGND VGND VPWR VPWR _06273_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_129_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10927_ _02522_ _02536_ VGND VGND VPWR VPWR _03226_ sky130_fd_sc_hd__and2_1
XFILLER_0_74_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13646_ _06013_ _06015_ VGND VGND VPWR VPWR _06198_ sky130_fd_sc_hd__or2_1
XFILLER_0_129_759 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10850__A2 _01410_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10858_ _03140_ _03139_ VGND VGND VPWR VPWR _03150_ sky130_fd_sc_hd__and2b_1
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13577_ _01249_ _02855_ _03785_ _02857_ VGND VGND VPWR VPWR _06122_ sky130_fd_sc_hd__and4_1
X_10789_ _00628_ _00650_ net54 _02312_ VGND VGND VPWR VPWR _03074_ sky130_fd_sc_hd__and4_1
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12528_ _04868_ _04985_ VGND VGND VPWR VPWR _04986_ sky130_fd_sc_hd__nand2_1
XFILLER_0_136_291 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12459_ _04898_ _04909_ VGND VGND VPWR VPWR _04910_ sky130_fd_sc_hd__or2_1
XFILLER_0_124_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14129_ _06649_ _06683_ _06725_ VGND VGND VPWR VPWR _06727_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_10_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10669__A2 _01411_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09670_ _01724_ _01726_ _01846_ VGND VGND VPWR VPWR _01847_ sky130_fd_sc_hd__o21a_1
XANTENNA__09381__A _01508_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08621_ _00698_ _00688_ VGND VGND VPWR VPWR _00700_ sky130_fd_sc_hd__and2b_1
XFILLER_0_77_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08552_ _00609_ _00610_ _00623_ VGND VGND VPWR VPWR _00624_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07503_ _01744_ _00311_ _04862_ _04873_ VGND VGND VPWR VPWR _04884_ sky130_fd_sc_hd__nand4_2
X_08483_ _00254_ _00328_ _00342_ VGND VGND VPWR VPWR _00549_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_76_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07434_ _03587_ _04015_ _04103_ _03576_ VGND VGND VPWR VPWR _04125_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10974__B _04939_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07365_ _00825_ _02773_ _02762_ VGND VGND VPWR VPWR _03367_ sky130_fd_sc_hd__a21o_1
XFILLER_0_128_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11789__C net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09104_ _01187_ _01227_ VGND VGND VPWR VPWR _01228_ sky130_fd_sc_hd__xor2_1
XFILLER_0_17_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07296_ _02499_ _02510_ _02587_ VGND VGND VPWR VPWR _02609_ sky130_fd_sc_hd__nand3_1
XFILLER_0_26_790 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09035_ _01117_ _01118_ _01151_ VGND VGND VPWR VPWR _01152_ sky130_fd_sc_hd__o21a_1
XFILLER_0_103_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07470__A1 _01197_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07470__B2 _04510_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09937_ _02136_ _02139_ VGND VGND VPWR VPWR _02140_ sky130_fd_sc_hd__and2_1
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09868_ _06873_ _00755_ _01260_ _06875_ VGND VGND VPWR VPWR _02064_ sky130_fd_sc_hd__a22o_1
X_08819_ _00741_ VGND VGND VPWR VPWR _00916_ sky130_fd_sc_hd__clkbuf_4
X_09799_ _01987_ _01988_ VGND VGND VPWR VPWR _01989_ sky130_fd_sc_hd__nor2_1
XTAP_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11609__A1 _00654_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11830_ _04217_ _04167_ VGND VGND VPWR VPWR _04218_ sky130_fd_sc_hd__nor2_1
XANTENNA__11609__B2 _00543_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11761_ _04122_ _04141_ VGND VGND VPWR VPWR _04142_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_68_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13500_ _06035_ _06036_ _01415_ _03680_ VGND VGND VPWR VPWR _06037_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_95_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10712_ _02959_ _02987_ _02988_ VGND VGND VPWR VPWR _02989_ sky130_fd_sc_hd__o21a_1
XFILLER_0_67_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11692_ _03510_ _01211_ _04063_ _04064_ VGND VGND VPWR VPWR _04066_ sky130_fd_sc_hd__o2bb2a_1
XTAP_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13431_ _05647_ _05663_ _05961_ VGND VGND VPWR VPWR _05962_ sky130_fd_sc_hd__and3_2
X_10643_ _02903_ _02912_ VGND VGND VPWR VPWR _02913_ sky130_fd_sc_hd__nand2_1
XANTENNA__12585__A2 _02158_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13362_ _05884_ _05885_ VGND VGND VPWR VPWR _05886_ sky130_fd_sc_hd__or2b_1
XFILLER_0_118_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10574_ _02824_ _02836_ VGND VGND VPWR VPWR _02837_ sky130_fd_sc_hd__nand2_1
Xrebuffer8 _04675_ VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12313_ _00459_ _01601_ _04747_ _04748_ _01288_ VGND VGND VPWR VPWR _04749_ sky130_fd_sc_hd__a32o_1
XFILLER_0_106_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13293_ _05801_ _05814_ VGND VGND VPWR VPWR _05815_ sky130_fd_sc_hd__nand2_1
XANTENNA__09738__B1 net52 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10108__C _05577_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12244_ _04671_ _04672_ VGND VGND VPWR VPWR _04673_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12175_ _03728_ _04017_ _04021_ _03725_ VGND VGND VPWR VPWR _04597_ sky130_fd_sc_hd__a211oi_1
X_11126_ _03443_ _03369_ VGND VGND VPWR VPWR _03445_ sky130_fd_sc_hd__or2_1
XANTENNA__10221__A1_N _02029_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11057_ _03365_ _03368_ VGND VGND VPWR VPWR _03369_ sky130_fd_sc_hd__and2_1
XANTENNA__09913__B _02040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10008_ _02211_ _02217_ VGND VGND VPWR VPWR _02218_ sky130_fd_sc_hd__nor2_1
XFILLER_0_64_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07433__B _03587_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07152__C net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11959_ _06417_ _02134_ _04359_ VGND VGND VPWR VPWR _04360_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_129_523 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10823__A2 net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_532 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13629_ _06074_ _06075_ _06178_ VGND VGND VPWR VPWR _06179_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_117_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08264__B _00298_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07150_ _00442_ _00989_ _01000_ _00901_ VGND VGND VPWR VPWR _01011_ sky130_fd_sc_hd__and4_1
XFILLER_0_54_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10587__A1 _00145_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10960__D _02189_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11000__A2 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07983_ _00020_ _00025_ VGND VGND VPWR VPWR _00027_ sky130_fd_sc_hd__and2_1
XANTENNA__13828__A2 _03680_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09722_ _01890_ _01903_ VGND VGND VPWR VPWR _01904_ sky130_fd_sc_hd__and2_1
XANTENNA__11839__A1 _03070_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11839__B2 _02456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09823__B _06820_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07624__A _05445_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12500__A2 _03696_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09653_ _01759_ _01760_ _01828_ VGND VGND VPWR VPWR _01829_ sky130_fd_sc_hd__or3b_2
XANTENNA__11791__D net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08604_ _00678_ _00680_ VGND VGND VPWR VPWR _00681_ sky130_fd_sc_hd__nor2_1
XANTENNA__10688__C net50 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09584_ _01486_ _01752_ VGND VGND VPWR VPWR _01753_ sky130_fd_sc_hd__or2b_1
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08535_ _00604_ VGND VGND VPWR VPWR _00605_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__08468__B1 _06875_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08466_ _03543_ _00095_ _00331_ _00330_ VGND VGND VPWR VPWR _00531_ sky130_fd_sc_hd__a31o_1
XFILLER_0_65_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07417_ net11 VGND VGND VPWR VPWR _03938_ sky130_fd_sc_hd__clkbuf_4
X_08397_ _00451_ _00452_ _04312_ VGND VGND VPWR VPWR _00455_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_80_619 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07348_ _03158_ _03169_ VGND VGND VPWR VPWR _03180_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_524 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07279_ _02248_ _02401_ _02412_ VGND VGND VPWR VPWR _02423_ sky130_fd_sc_hd__a21o_2
XFILLER_0_60_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09286__A _01309_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09018_ _03543_ _00144_ _00994_ _00993_ VGND VGND VPWR VPWR _01134_ sky130_fd_sc_hd__a31o_1
XFILLER_0_131_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10290_ _02156_ _02524_ _02525_ VGND VGND VPWR VPWR _02526_ sky130_fd_sc_hd__a21bo_1
XANTENNA__11527__B1 _03690_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13819__A2 _01955_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13536__A _02722_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13980_ _06157_ _06564_ VGND VGND VPWR VPWR _06565_ sky130_fd_sc_hd__or2_1
X_12931_ _04536_ _05428_ VGND VGND VPWR VPWR _05429_ sky130_fd_sc_hd__xnor2_4
XANTENNA__07534__A _01361_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13255__B _05546_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12862_ _05337_ _05352_ VGND VGND VPWR VPWR _05353_ sky130_fd_sc_hd__xor2_2
XTAP_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11813_ _04194_ _04195_ _04198_ VGND VGND VPWR VPWR _04199_ sky130_fd_sc_hd__o21a_1
XTAP_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12793_ _02728_ _05100_ _05276_ VGND VGND VPWR VPWR _05277_ sky130_fd_sc_hd__a21bo_1
XTAP_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11744_ _04120_ _04117_ VGND VGND VPWR VPWR _04123_ sky130_fd_sc_hd__nand2_1
XFILLER_0_139_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07682__A1 _01076_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11675_ _04041_ _04046_ VGND VGND VPWR VPWR _04047_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10018__B1 _00379_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13414_ _05898_ _05942_ VGND VGND VPWR VPWR _05943_ sky130_fd_sc_hd__nand2_1
X_10626_ _02842_ _02893_ VGND VGND VPWR VPWR _02895_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10569__A1 _00819_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09423__A2 _00745_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_855 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07434__A1 _03587_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13345_ _05865_ _05866_ VGND VGND VPWR VPWR _05867_ sky130_fd_sc_hd__nor2_1
XANTENNA__07434__B2 _03576_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10557_ _02803_ _02802_ VGND VGND VPWR VPWR _02819_ sky130_fd_sc_hd__and2b_1
XFILLER_0_59_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13276_ _05472_ _05799_ VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__xor2_4
X_10488_ _02736_ VGND VGND VPWR VPWR _02743_ sky130_fd_sc_hd__clkbuf_4
X_12227_ _01517_ _03738_ _03744_ _01518_ VGND VGND VPWR VPWR _04655_ sky130_fd_sc_hd__a22o_1
XANTENNA__07737__A2 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12158_ _04570_ _04571_ VGND VGND VPWR VPWR _04579_ sky130_fd_sc_hd__nand2_1
X_11109_ _03409_ _03425_ VGND VGND VPWR VPWR _03426_ sky130_fd_sc_hd__nand2_1
X_12089_ _04500_ _04502_ VGND VGND VPWR VPWR _04503_ sky130_fd_sc_hd__xor2_2
XANTENNA__10789__B _00650_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07444__A _01372_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08259__B _00138_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08320_ _00352_ _00369_ _00370_ VGND VGND VPWR VPWR _00371_ sky130_fd_sc_hd__o21ai_2
XANTENNA__12797__A2 _01933_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08251_ _06428_ _06450_ _00293_ _00294_ VGND VGND VPWR VPWR _00295_ sky130_fd_sc_hd__and4_1
XFILLER_0_46_159 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07202_ _01230_ _00300_ VGND VGND VPWR VPWR _01580_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08182_ _03488_ _03609_ _00225_ VGND VGND VPWR VPWR _00226_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_27_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_518 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07133_ _00694_ _00814_ VGND VGND VPWR VPWR _00825_ sky130_fd_sc_hd__nor2_1
XFILLER_0_70_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09818__B _01260_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07966_ _01076_ _07010_ net38 _01120_ VGND VGND VPWR VPWR _00010_ sky130_fd_sc_hd__a22o_1
XANTENNA__12260__A _00376_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09705_ _01883_ _01884_ VGND VGND VPWR VPWR _01885_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07897_ _07024_ _07025_ VGND VGND VPWR VPWR _07026_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09636_ _01177_ _01808_ _01809_ VGND VGND VPWR VPWR _01811_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_69_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13803__B _03679_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09567_ _01476_ _01734_ VGND VGND VPWR VPWR _01735_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08518_ _00580_ _00586_ VGND VGND VPWR VPWR _00587_ sky130_fd_sc_hd__xor2_2
XFILLER_0_38_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09498_ _01657_ _01658_ VGND VGND VPWR VPWR _01659_ sky130_fd_sc_hd__xor2_1
XFILLER_0_92_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08449_ _00316_ _00511_ VGND VGND VPWR VPWR _00512_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11460_ _03808_ _03810_ VGND VGND VPWR VPWR _03811_ sky130_fd_sc_hd__or2b_1
XFILLER_0_18_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07416__A1 _00311_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10411_ _02657_ _02658_ VGND VGND VPWR VPWR _02659_ sky130_fd_sc_hd__nand2_1
X_11391_ _03733_ _03734_ VGND VGND VPWR VPWR _03735_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13130_ _05631_ _05647_ VGND VGND VPWR VPWR _05648_ sky130_fd_sc_hd__and2_4
X_10342_ _02542_ _02582_ VGND VGND VPWR VPWR _02583_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_104_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13061_ _05559_ _05571_ VGND VGND VPWR VPWR _05572_ sky130_fd_sc_hd__xnor2_2
X_10273_ _03576_ _00989_ _02312_ VGND VGND VPWR VPWR _02507_ sky130_fd_sc_hd__and3_1
X_12012_ _04416_ _04417_ VGND VGND VPWR VPWR _04418_ sky130_fd_sc_hd__nor2_1
XANTENNA__07264__A _02116_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13963_ _06544_ _06545_ VGND VGND VPWR VPWR _06546_ sky130_fd_sc_hd__nor2_1
XANTENNA__08079__B _06964_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12914_ _05259_ _05305_ VGND VGND VPWR VPWR _05410_ sky130_fd_sc_hd__nand2_1
X_13894_ _06468_ _06469_ VGND VGND VPWR VPWR _06470_ sky130_fd_sc_hd__or2b_1
XFILLER_0_88_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12845_ _05286_ _05333_ VGND VGND VPWR VPWR _05334_ sky130_fd_sc_hd__or2_1
XTAP_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14097__A _06684_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12776_ _05256_ _05257_ VGND VGND VPWR VPWR _05259_ sky130_fd_sc_hd__xor2_2
XTAP_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08095__A _00138_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11727_ _04102_ _04104_ VGND VGND VPWR VPWR _04105_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12217__A1_N _00458_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_142_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11658_ _03862_ _04008_ VGND VGND VPWR VPWR _04029_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_83_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09919__A _01960_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11739__B1 _01289_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10609_ _02873_ _02875_ VGND VGND VPWR VPWR _02876_ sky130_fd_sc_hd__nand2_1
XFILLER_0_142_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11589_ _01155_ _01957_ _03952_ VGND VGND VPWR VPWR _03953_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_40_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_140 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12345__A _00915_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07439__A net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13328_ _05843_ _05849_ VGND VGND VPWR VPWR _05850_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08261__C _02018_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13259_ _05596_ _05545_ _05783_ VGND VGND VPWR VPWR _05784_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_20_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07820_ _06862_ _06948_ VGND VGND VPWR VPWR _06949_ sky130_fd_sc_hd__nor2_1
XANTENNA__12080__A _02246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07751_ _06878_ _06879_ VGND VGND VPWR VPWR _06880_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_79_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10478__B1 _02731_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07682_ _01076_ _03499_ _06797_ _06802_ VGND VGND VPWR VPWR _06809_ sky130_fd_sc_hd__a31o_1
XFILLER_0_79_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09421_ _00138_ _00742_ VGND VGND VPWR VPWR _01575_ sky130_fd_sc_hd__nand2_1
XANTENNA__11690__A2 _00571_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09352_ _01364_ _01497_ VGND VGND VPWR VPWR _01499_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09635__A2 _01177_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08303_ _03839_ _00351_ VGND VGND VPWR VPWR _00352_ sky130_fd_sc_hd__and2_2
XFILLER_0_75_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09283_ _01360_ _01422_ VGND VGND VPWR VPWR _01424_ sky130_fd_sc_hd__nor2_1
XANTENNA__07340__C _02105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11442__A2 _02133_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08234_ _00273_ _00276_ VGND VGND VPWR VPWR _00278_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_682 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08165_ _06845_ _06846_ VGND VGND VPWR VPWR _00209_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07116_ net28 VGND VGND VPWR VPWR _00639_ sky130_fd_sc_hd__buf_8
XANTENNA__12942__A2 _02150_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08096_ _02018_ _04895_ _04928_ _05478_ VGND VGND VPWR VPWR _00140_ sky130_fd_sc_hd__a22o_1
XFILLER_0_113_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08998_ _01057_ _01111_ VGND VGND VPWR VPWR _01112_ sky130_fd_sc_hd__xnor2_2
XANTENNA__10503__A _02758_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07949_ _07037_ _07076_ VGND VGND VPWR VPWR _07078_ sky130_fd_sc_hd__nor2_1
XANTENNA__10222__B _01564_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10960_ _00145_ _00310_ _02187_ _02189_ VGND VGND VPWR VPWR _03262_ sky130_fd_sc_hd__and4_1
XANTENNA__07334__B1 _03015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09619_ _01261_ _01576_ _01579_ VGND VGND VPWR VPWR _01792_ sky130_fd_sc_hd__and3_1
X_10891_ _03176_ _03184_ _03185_ VGND VGND VPWR VPWR _03186_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_85_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12630_ _05096_ _05086_ VGND VGND VPWR VPWR _05098_ sky130_fd_sc_hd__or2_1
XANTENNA__09087__B1 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12561_ _00390_ _01066_ _05020_ VGND VGND VPWR VPWR _05022_ sky130_fd_sc_hd__and3_1
XFILLER_0_66_777 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11512_ _03865_ _03867_ VGND VGND VPWR VPWR _03868_ sky130_fd_sc_hd__nand2_1
XANTENNA__09739__A _04169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12492_ _00780_ _00777_ _03685_ _00423_ VGND VGND VPWR VPWR _04946_ sky130_fd_sc_hd__and4_1
XFILLER_0_135_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14231_ _00249_ _00361_ VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__xnor2_1
XFILLER_0_124_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11443_ _06964_ _00121_ _02133_ _02459_ VGND VGND VPWR VPWR _03792_ sky130_fd_sc_hd__and4_1
XFILLER_0_22_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12394__B1 _00571_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14162_ _06730_ _06731_ _06732_ VGND VGND VPWR VPWR _06761_ sky130_fd_sc_hd__and3_1
XFILLER_0_33_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08062__A1 _06472_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11374_ _01312_ _00544_ _01957_ _03690_ VGND VGND VPWR VPWR _03716_ sky130_fd_sc_hd__and4_2
XFILLER_0_104_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13113_ _04601_ _04628_ VGND VGND VPWR VPWR _05629_ sky130_fd_sc_hd__xor2_1
X_10325_ _04862_ net4 _00780_ VGND VGND VPWR VPWR _02564_ sky130_fd_sc_hd__and3_1
X_14093_ _06686_ _05848_ VGND VGND VPWR VPWR _06688_ sky130_fd_sc_hd__or2b_1
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13044_ _04573_ _05552_ VGND VGND VPWR VPWR _05553_ sky130_fd_sc_hd__nand2_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10256_ _02487_ _02488_ VGND VGND VPWR VPWR _02490_ sky130_fd_sc_hd__or2_2
XANTENNA__13708__B _02759_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07706__B net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10187_ _03499_ _06821_ net13 _00730_ VGND VGND VPWR VPWR _02414_ sky130_fd_sc_hd__and4_1
X_13946_ _06511_ _06513_ VGND VGND VPWR VPWR _06528_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08818__A _00914_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13877_ _06445_ _06449_ _06436_ VGND VGND VPWR VPWR _06452_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07441__B _04169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12828_ _04601_ _04628_ _05315_ VGND VGND VPWR VPWR _05316_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_29_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12759_ _00457_ _03744_ VGND VGND VPWR VPWR _05240_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12385__B1 _00734_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07169__A _00880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09970_ _02171_ _01060_ _01413_ _02259_ VGND VGND VPWR VPWR _02176_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_110_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08921_ _00833_ _01026_ _01025_ VGND VGND VPWR VPWR _01028_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08852_ _00950_ _00951_ VGND VGND VPWR VPWR _00952_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11419__A _06775_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07803_ _06929_ _06931_ VGND VGND VPWR VPWR _06932_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_137_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08783_ _00874_ _00876_ VGND VGND VPWR VPWR _00877_ sky130_fd_sc_hd__xnor2_2
XANTENNA__07335__C _00355_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07734_ _06852_ _06861_ VGND VGND VPWR VPWR _06863_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10977__B _00607_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07665_ _06626_ _06637_ _06208_ VGND VGND VPWR VPWR _06648_ sky130_fd_sc_hd__and3_1
XANTENNA__08795__B1_N _00598_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11663__A2 _00414_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09404_ _01500_ _01555_ VGND VGND VPWR VPWR _01556_ sky130_fd_sc_hd__xnor2_1
X_07596_ _05868_ _05879_ VGND VGND VPWR VPWR _05890_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09335_ _01346_ VGND VGND VPWR VPWR _01480_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09266_ _01403_ _01404_ VGND VGND VPWR VPWR _01406_ sky130_fd_sc_hd__xor2_1
XFILLER_0_90_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08463__A _00519_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_142 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08217_ _00125_ _00124_ VGND VGND VPWR VPWR _00261_ sky130_fd_sc_hd__and2b_1
XFILLER_0_62_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09197_ _01005_ _01146_ VGND VGND VPWR VPWR _01330_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08148_ _05346_ VGND VGND VPWR VPWR _00192_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08595__A2 _00257_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13809__A _02187_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08079_ _05566_ _06964_ _00122_ VGND VGND VPWR VPWR _00123_ sky130_fd_sc_hd__and3_1
XFILLER_0_30_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10110_ _02177_ _02328_ VGND VGND VPWR VPWR _02329_ sky130_fd_sc_hd__and2_1
X_11090_ _02558_ _03327_ VGND VGND VPWR VPWR _03405_ sky130_fd_sc_hd__and2_1
XFILLER_0_101_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10041_ _01841_ _01844_ _02252_ VGND VGND VPWR VPWR _02254_ sky130_fd_sc_hd__nor3_1
XANTENNA__11351__A1 _00544_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11351__B2 _03690_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13800_ _02187_ _03682_ VGND VGND VPWR VPWR _06367_ sky130_fd_sc_hd__nand2_1
XANTENNA__09741__B net50 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11992_ _04394_ _04395_ VGND VGND VPWR VPWR _04396_ sky130_fd_sc_hd__nand2_2
XANTENNA__07542__A _00333_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10943_ _03073_ _03100_ VGND VGND VPWR VPWR _03243_ sky130_fd_sc_hd__and2_1
XFILLER_0_86_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13731_ _06286_ _06284_ VGND VGND VPWR VPWR _06291_ sky130_fd_sc_hd__and2b_1
XFILLER_0_98_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13662_ _06207_ _06209_ _06211_ VGND VGND VPWR VPWR _06215_ sky130_fd_sc_hd__nand3_1
XFILLER_0_42_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10874_ _03145_ _03148_ _03166_ _03142_ VGND VGND VPWR VPWR _03167_ sky130_fd_sc_hd__a211o_1
XFILLER_0_78_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12613_ _05068_ _05069_ VGND VGND VPWR VPWR _05079_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_66_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13593_ _06136_ _06138_ VGND VGND VPWR VPWR _06139_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_120 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09469__A _01626_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12544_ _04996_ _05002_ VGND VGND VPWR VPWR _05003_ sky130_fd_sc_hd__or2b_1
XFILLER_0_81_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12475_ _04924_ _04921_ VGND VGND VPWR VPWR _04927_ sky130_fd_sc_hd__and2b_1
XFILLER_0_41_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14214_ net157 _02423_ VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__xor2_4
X_11426_ _03760_ _03761_ VGND VGND VPWR VPWR _03774_ sky130_fd_sc_hd__xor2_1
XFILLER_0_1_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14145_ _06714_ _06742_ VGND VGND VPWR VPWR _06743_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11357_ _01312_ _03697_ _03693_ _03694_ VGND VGND VPWR VPWR _03698_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_22_688 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08820__B _00159_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10308_ _02350_ _02352_ VGND VGND VPWR VPWR _02546_ sky130_fd_sc_hd__nand2_1
X_14076_ _06074_ _04013_ _06667_ VGND VGND VPWR VPWR _06670_ sky130_fd_sc_hd__a21oi_1
XTAP_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output79_A net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11288_ _03484_ _03486_ VGND VGND VPWR VPWR _03623_ sky130_fd_sc_hd__xor2_4
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13027_ _02480_ _04577_ _04579_ _05534_ VGND VGND VPWR VPWR _05535_ sky130_fd_sc_hd__a31o_1
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10239_ _02439_ _02470_ VGND VGND VPWR VPWR _02471_ sky130_fd_sc_hd__xor2_2
XANTENNA__09932__A _02133_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xrebuffer18 _04400_ VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__clkbuf_1
Xrebuffer29 _00716_ VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__buf_1
XFILLER_0_16_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13929_ _06220_ _06508_ VGND VGND VPWR VPWR _06509_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_76_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07450_ _04246_ _04290_ VGND VGND VPWR VPWR _04301_ sky130_fd_sc_hd__xnor2_1
X_07381_ _03532_ VGND VGND VPWR VPWR _03543_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_72_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09120_ _01231_ _01244_ VGND VGND VPWR VPWR _01245_ sky130_fd_sc_hd__nand2_1
XANTENNA__09471__B1 _01309_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08283__A _00377_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_235 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09051_ _00987_ _01168_ _01169_ VGND VGND VPWR VPWR _01170_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_5_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08002_ _00043_ _00045_ VGND VGND VPWR VPWR _00046_ sky130_fd_sc_hd__and2_1
XFILLER_0_115_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09953_ _04268_ _01546_ _02156_ _01372_ VGND VGND VPWR VPWR _02157_ sky130_fd_sc_hd__a22o_1
XANTENNA__12252__B _02120_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08904_ _00388_ _00112_ _00114_ _03004_ VGND VGND VPWR VPWR _01009_ sky130_fd_sc_hd__a22oi_1
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09884_ _02076_ _02080_ VGND VGND VPWR VPWR _02081_ sky130_fd_sc_hd__xor2_1
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08835_ _00917_ _00744_ _00918_ _00931_ VGND VGND VPWR VPWR _00933_ sky130_fd_sc_hd__o31ai_2
X_08766_ _00310_ VGND VGND VPWR VPWR _00859_ sky130_fd_sc_hd__clkbuf_4
X_07717_ _06836_ _06838_ VGND VGND VPWR VPWR _06846_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_68_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08697_ _00782_ VGND VGND VPWR VPWR _00783_ sky130_fd_sc_hd__buf_2
X_07648_ _05588_ VGND VGND VPWR VPWR _06461_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_95_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13389__A2 _02673_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07579_ _05654_ _05698_ _05665_ VGND VGND VPWR VPWR _05720_ sky130_fd_sc_hd__and3_1
X_09318_ _01337_ _01342_ _01460_ VGND VGND VPWR VPWR _01462_ sky130_fd_sc_hd__o21a_1
XANTENNA__12597__B1 _02849_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10590_ _02306_ VGND VGND VPWR VPWR _02855_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_90_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09249_ _01382_ _01386_ VGND VGND VPWR VPWR _01387_ sky130_fd_sc_hd__xor2_1
XFILLER_0_8_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10228__A net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12260_ _00376_ _00378_ _01180_ _01249_ VGND VGND VPWR VPWR _04691_ sky130_fd_sc_hd__and4_2
XFILLER_0_105_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11211_ _02502_ _02541_ _02582_ VGND VGND VPWR VPWR _03538_ sky130_fd_sc_hd__a21oi_2
X_12191_ _03533_ _03514_ VGND VGND VPWR VPWR _04615_ sky130_fd_sc_hd__or2b_1
XANTENNA__10375__A2 _00413_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11142_ _03250_ _03449_ VGND VGND VPWR VPWR _03462_ sky130_fd_sc_hd__xor2_2
XFILLER_0_101_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput65 net65 VGND VGND VPWR VPWR prod[0] sky130_fd_sc_hd__clkbuf_4
Xoutput76 net76 VGND VGND VPWR VPWR prod[1] sky130_fd_sc_hd__clkbuf_4
Xoutput87 net87 VGND VGND VPWR VPWR prod[2] sky130_fd_sc_hd__buf_2
X_11073_ _03384_ _03385_ VGND VGND VPWR VPWR _03386_ sky130_fd_sc_hd__nor2_1
Xoutput98 net98 VGND VGND VPWR VPWR prod[3] sky130_fd_sc_hd__clkbuf_4
X_10024_ _02233_ _02234_ VGND VGND VPWR VPWR _02235_ sky130_fd_sc_hd__nand2_2
XANTENNA__08368__A net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11975_ _04374_ _04376_ VGND VGND VPWR VPWR _04377_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output117_A net117 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13714_ _02426_ _02759_ _06271_ VGND VGND VPWR VPWR _06272_ sky130_fd_sc_hd__and3_1
X_10926_ _02467_ _02758_ VGND VGND VPWR VPWR _03225_ sky130_fd_sc_hd__and2_1
XFILLER_0_128_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13645_ _06193_ _06194_ VGND VGND VPWR VPWR _06196_ sky130_fd_sc_hd__nor2_1
X_10857_ _05588_ _01410_ _02525_ _02524_ _02304_ VGND VGND VPWR VPWR _03149_ sky130_fd_sc_hd__a32o_1
XFILLER_0_67_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10788_ _03063_ _03071_ VGND VGND VPWR VPWR _03073_ sky130_fd_sc_hd__xor2_1
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13576_ _02855_ _03785_ VGND VGND VPWR VPWR _06121_ sky130_fd_sc_hd__nand2_1
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12527_ _04866_ _04867_ VGND VGND VPWR VPWR _04985_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12458_ _04905_ _04907_ _04908_ VGND VGND VPWR VPWR _04909_ sky130_fd_sc_hd__a21o_1
XFILLER_0_112_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11409_ _03752_ _03753_ _03749_ VGND VGND VPWR VPWR _03755_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12389_ _00779_ _01586_ _01584_ _00784_ VGND VGND VPWR VPWR _04833_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__07447__A _01230_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14128_ _06649_ _06683_ _06725_ VGND VGND VPWR VPWR _06726_ sky130_fd_sc_hd__or3b_2
XFILLER_0_10_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14059_ _06062_ _06093_ _06061_ VGND VGND VPWR VPWR _06651_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_118_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08620_ _00688_ _00698_ VGND VGND VPWR VPWR _00699_ sky130_fd_sc_hd__and2b_1
XANTENNA__07182__A _01295_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08551_ _00621_ _00622_ VGND VGND VPWR VPWR _00623_ sky130_fd_sc_hd__xor2_1
X_07502_ net4 VGND VGND VPWR VPWR _04873_ sky130_fd_sc_hd__buf_4
XFILLER_0_134_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08482_ _00525_ _00547_ VGND VGND VPWR VPWR _00548_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07433_ _03576_ _03587_ _04015_ _04103_ VGND VGND VPWR VPWR _04114_ sky130_fd_sc_hd__and4_1
XANTENNA__10974__C _00460_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12579__B1 _02720_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07364_ _03334_ _03345_ VGND VGND VPWR VPWR _03356_ sky130_fd_sc_hd__or2b_1
XFILLER_0_18_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09103_ _01189_ _01226_ VGND VGND VPWR VPWR _01227_ sky130_fd_sc_hd__xor2_2
XANTENNA__11789__D net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07295_ _02499_ _02510_ _02587_ VGND VGND VPWR VPWR _02598_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_72_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09034_ _01149_ _01150_ VGND VGND VPWR VPWR _01151_ sky130_fd_sc_hd__nand2_1
XFILLER_0_143_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07470__A2 _04367_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08460__B _00523_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09936_ _02137_ VGND VGND VPWR VPWR _02139_ sky130_fd_sc_hd__inv_2
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09867_ _03521_ _01260_ _02016_ _02015_ VGND VGND VPWR VPWR _02063_ sky130_fd_sc_hd__a31o_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07804__B _05291_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08818_ _00914_ VGND VGND VPWR VPWR _00915_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09798_ _03059_ _01585_ _01983_ _01986_ VGND VGND VPWR VPWR _01988_ sky130_fd_sc_hd__and4_1
XANTENNA__07092__A _00366_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07930__B1 net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08749_ _00664_ _00838_ VGND VGND VPWR VPWR _00840_ sky130_fd_sc_hd__or2_1
XANTENNA__11609__A2 _01181_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11760_ _04134_ _04137_ _04139_ _04140_ VGND VGND VPWR VPWR _04141_ sky130_fd_sc_hd__a31o_1
XTAP_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10293__A1 _05577_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10711_ _02945_ _02947_ VGND VGND VPWR VPWR _02988_ sky130_fd_sc_hd__xor2_1
XTAP_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11691_ _04063_ _04064_ _03510_ _01211_ VGND VGND VPWR VPWR _04065_ sky130_fd_sc_hd__and4bb_1
XTAP_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11342__A _02459_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10642_ _02910_ _02911_ VGND VGND VPWR VPWR _02912_ sky130_fd_sc_hd__nor2_1
X_13430_ _05424_ _05631_ VGND VGND VPWR VPWR _05961_ sky130_fd_sc_hd__and2b_1
XFILLER_0_119_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13361_ _05337_ _05352_ _05883_ VGND VGND VPWR VPWR _05885_ sky130_fd_sc_hd__nand3_1
XFILLER_0_106_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10573_ _02821_ _02823_ VGND VGND VPWR VPWR _02836_ sky130_fd_sc_hd__or2_1
XFILLER_0_51_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12312_ _00415_ _00607_ _01664_ VGND VGND VPWR VPWR _04748_ sky130_fd_sc_hd__and3_1
Xrebuffer9 _05037_ VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__buf_1
X_13292_ _05712_ _05725_ VGND VGND VPWR VPWR _05814_ sky130_fd_sc_hd__and2_1
XANTENNA__09738__A1 _00891_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12243_ _04665_ _04668_ _04670_ VGND VGND VPWR VPWR _04672_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09738__B2 _03587_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12742__B1 _02134_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12174_ _04025_ _04028_ _04032_ _04595_ VGND VGND VPWR VPWR _04596_ sky130_fd_sc_hd__or4b_4
XFILLER_0_31_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11125_ _03298_ _03442_ VGND VGND VPWR VPWR _03443_ sky130_fd_sc_hd__nor2_1
X_11056_ _03289_ _03366_ VGND VGND VPWR VPWR _03368_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09913__C _01179_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10007_ _02212_ _02216_ VGND VGND VPWR VPWR _02217_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09910__A1 _00333_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10421__A _02127_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08098__A _05027_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07433__C _04015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07152__D net61 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11958_ _00138_ _02459_ VGND VGND VPWR VPWR _04359_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10909_ _03199_ _03203_ VGND VGND VPWR VPWR _03206_ sky130_fd_sc_hd__nor2_1
XFILLER_0_80_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11889_ _04104_ _04040_ VGND VGND VPWR VPWR _04283_ sky130_fd_sc_hd__and2b_1
X_13628_ _06176_ _06169_ _06173_ VGND VGND VPWR VPWR _06178_ sky130_fd_sc_hd__and3_1
XFILLER_0_27_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13559_ _06071_ _06101_ VGND VGND VPWR VPWR _06102_ sky130_fd_sc_hd__and2_1
XANTENNA__10587__A2 _01413_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07177__A _01208_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07982_ _00020_ _00025_ VGND VGND VPWR VPWR _00026_ sky130_fd_sc_hd__nor2_1
X_09721_ _01677_ _01902_ VGND VGND VPWR VPWR _01903_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11839__A2 _01955_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09823__C net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11427__A _00004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07624__B _05467_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09652_ _01825_ _01827_ VGND VGND VPWR VPWR _01828_ sky130_fd_sc_hd__xor2_4
XANTENNA__10331__A net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08603_ _00280_ _00482_ _00679_ VGND VGND VPWR VPWR _00680_ sky130_fd_sc_hd__a21oi_1
X_09583_ _01721_ _01751_ VGND VGND VPWR VPWR _01752_ sky130_fd_sc_hd__xor2_2
XFILLER_0_77_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08534_ net46 VGND VGND VPWR VPWR _00604_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_49_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08468__A1 _02993_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08468__B2 _05203_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10275__A1 net57 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08465_ _00335_ _00338_ VGND VGND VPWR VPWR _00529_ sky130_fd_sc_hd__and2b_1
XFILLER_0_77_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12258__A _00378_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07416_ _00311_ _03762_ _03806_ _03795_ VGND VGND VPWR VPWR _03927_ sky130_fd_sc_hd__a31o_1
XFILLER_0_135_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08396_ _04312_ _00451_ _00452_ VGND VGND VPWR VPWR _00454_ sky130_fd_sc_hd__and3_1
XFILLER_0_70_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07347_ _01044_ _03147_ _00880_ net26 VGND VGND VPWR VPWR _03169_ sky130_fd_sc_hd__nand4_1
XFILLER_0_18_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07278_ _02215_ _02237_ VGND VGND VPWR VPWR _02412_ sky130_fd_sc_hd__and2_1
X_09017_ _01018_ _01132_ VGND VGND VPWR VPWR _01133_ sky130_fd_sc_hd__xor2_1
XFILLER_0_115_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11527__A1 _01312_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11527__B2 _01155_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07087__A _00311_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12721__A _00391_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09919_ _01960_ VGND VGND VPWR VPWR _02120_ sky130_fd_sc_hd__clkbuf_4
X_12930_ _04491_ _05427_ VGND VGND VPWR VPWR _05428_ sky130_fd_sc_hd__nand2_2
XANTENNA__07534__B _05181_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12861_ _05350_ _05351_ VGND VGND VPWR VPWR _05352_ sky130_fd_sc_hd__and2_1
XTAP_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11812_ _04161_ _04197_ VGND VGND VPWR VPWR _04198_ sky130_fd_sc_hd__xor2_1
XTAP_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12792_ _00392_ _02723_ _02727_ _00389_ VGND VGND VPWR VPWR _05276_ sky130_fd_sc_hd__a22o_1
XTAP_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11743_ _04106_ _04121_ VGND VGND VPWR VPWR _04122_ sky130_fd_sc_hd__xnor2_2
XTAP_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07682__A2 _03499_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11674_ _04044_ _04045_ VGND VGND VPWR VPWR _04046_ sky130_fd_sc_hd__nor2_1
XFILLER_0_138_398 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10018__A1 _04939_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10018__B2 _04917_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13413_ _05406_ _05941_ VGND VGND VPWR VPWR _05942_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10625_ _02865_ _02892_ VGND VGND VPWR VPWR _02893_ sky130_fd_sc_hd__xor2_1
XANTENNA__10569__A2 _01934_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07434__A2 _04015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10556_ _02814_ _02816_ VGND VGND VPWR VPWR _02818_ sky130_fd_sc_hd__or2_1
X_13344_ _05854_ _05336_ _05864_ VGND VGND VPWR VPWR _05866_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_52_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13275_ _05795_ _05798_ VGND VGND VPWR VPWR _05799_ sky130_fd_sc_hd__nand2_2
X_10487_ _02737_ VGND VGND VPWR VPWR _02742_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_121_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12226_ _01518_ _01517_ _03738_ _03744_ VGND VGND VPWR VPWR _04654_ sky130_fd_sc_hd__nand4_2
XFILLER_0_121_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12157_ _04566_ _04574_ VGND VGND VPWR VPWR _04578_ sky130_fd_sc_hd__nor2_2
X_11108_ _03406_ _03408_ VGND VGND VPWR VPWR _03425_ sky130_fd_sc_hd__or2_1
X_12088_ _04353_ _04354_ _04355_ _04423_ _04501_ VGND VGND VPWR VPWR _04502_ sky130_fd_sc_hd__a41o_2
XANTENNA__10789__C net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11039_ _03347_ _03348_ VGND VGND VPWR VPWR _03349_ sky130_fd_sc_hd__xnor2_2
XANTENNA__07444__B _04026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08259__C _04906_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08250_ _00151_ VGND VGND VPWR VPWR _00294_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_86_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_398 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07201_ _01536_ _01558_ VGND VGND VPWR VPWR _01569_ sky130_fd_sc_hd__xor2_2
X_08181_ _03488_ _03609_ _03048_ VGND VGND VPWR VPWR _00225_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_15_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07132_ _00770_ _00803_ VGND VGND VPWR VPWR _00814_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11710__A _00258_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07965_ _01120_ net37 _07013_ _07012_ VGND VGND VPWR VPWR _00009_ sky130_fd_sc_hd__a31o_1
XANTENNA__12260__B _00378_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09704_ _00388_ _00459_ VGND VGND VPWR VPWR _01884_ sky130_fd_sc_hd__and2_1
X_07896_ _02719_ _03499_ VGND VGND VPWR VPWR _07025_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09635_ _01197_ _01177_ _01246_ _04510_ VGND VGND VPWR VPWR _01809_ sky130_fd_sc_hd__a22o_1
XFILLER_0_139_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09566_ _01731_ _01732_ VGND VGND VPWR VPWR _01734_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08517_ _00583_ _00585_ VGND VGND VPWR VPWR _00586_ sky130_fd_sc_hd__nor2_1
XANTENNA__13091__B _04627_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09497_ _04268_ net49 VGND VGND VPWR VPWR _01658_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08448_ _00509_ _00510_ VGND VGND VPWR VPWR _00511_ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08379_ _02335_ _00389_ VGND VGND VPWR VPWR _00435_ sky130_fd_sc_hd__and2_1
XFILLER_0_34_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10410_ _02652_ _02656_ VGND VGND VPWR VPWR _02658_ sky130_fd_sc_hd__or2_1
XFILLER_0_116_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11390_ _03732_ _03723_ VGND VGND VPWR VPWR _03734_ sky130_fd_sc_hd__and2b_1
XANTENNA__07416__A2 _03762_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10341_ _02579_ _02581_ VGND VGND VPWR VPWR _02582_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_103_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10420__A1 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13060_ _05549_ _05556_ VGND VGND VPWR VPWR _05571_ sky130_fd_sc_hd__xnor2_1
X_10272_ _02309_ _02310_ VGND VGND VPWR VPWR _02506_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12011_ _04337_ _04415_ VGND VGND VPWR VPWR _04417_ sky130_fd_sc_hd__nor2_1
XANTENNA__07545__A _02335_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13962_ _06541_ _06542_ VGND VGND VPWR VPWR _06545_ sky130_fd_sc_hd__nor2_1
X_12913_ _05362_ _05408_ VGND VGND VPWR VPWR _05409_ sky130_fd_sc_hd__xnor2_1
X_13893_ _05929_ _05936_ _05930_ VGND VGND VPWR VPWR _06469_ sky130_fd_sc_hd__a21bo_1
XTAP_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12844_ _05325_ _05332_ VGND VGND VPWR VPWR _05333_ sky130_fd_sc_hd__xor2_1
XFILLER_0_69_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12775_ _04712_ _04724_ _04711_ VGND VGND VPWR VPWR _05257_ sky130_fd_sc_hd__a21o_1
XFILLER_0_56_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08095__B _02007_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11726_ _04083_ _04101_ VGND VGND VPWR VPWR _04104_ sky130_fd_sc_hd__and2_1
XFILLER_0_28_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11657_ _04012_ _04027_ VGND VGND VPWR VPWR _04028_ sky130_fd_sc_hd__nand2_2
XFILLER_0_37_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11739__A1 _00654_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11739__B2 _00543_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10608_ _02869_ _02874_ VGND VGND VPWR VPWR _02875_ sky130_fd_sc_hd__xnor2_1
X_11588_ _03950_ _03943_ _03947_ VGND VGND VPWR VPWR _03952_ sky130_fd_sc_hd__and3_1
XANTENNA__12345__B _01664_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13327_ _05820_ _05842_ _05848_ VGND VGND VPWR VPWR _05849_ sky130_fd_sc_hd__o21ba_1
X_10539_ _02797_ _02798_ VGND VGND VPWR VPWR _02799_ sky130_fd_sc_hd__or2b_1
XFILLER_0_24_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08261__D _00143_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09935__A _02127_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13258_ _05519_ _05523_ VGND VGND VPWR VPWR _05783_ sky130_fd_sc_hd__and2_1
XFILLER_0_122_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12209_ _00379_ _03682_ _04634_ _04630_ VGND VGND VPWR VPWR _04635_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__10175__B1 _03718_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13189_ _05694_ _05712_ VGND VGND VPWR VPWR _05713_ sky130_fd_sc_hd__nand2_1
XANTENNA__12080__B _02426_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07750_ _06829_ _06849_ _06827_ VGND VGND VPWR VPWR _06879_ sky130_fd_sc_hd__a21oi_2
XANTENNA__09868__B1 _01260_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10478__A1 _01472_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07681_ net1 net12 net35 net34 VGND VGND VPWR VPWR _06802_ sky130_fd_sc_hd__and4_1
XANTENNA__10478__B2 _00636_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13192__A _05464_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09420_ _01193_ _01199_ _01265_ VGND VGND VPWR VPWR _01574_ sky130_fd_sc_hd__and3_1
XANTENNA__08286__A _03532_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09351_ _01364_ _01497_ VGND VGND VPWR VPWR _01498_ sky130_fd_sc_hd__and2_1
XFILLER_0_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08302_ _03751_ _03828_ VGND VGND VPWR VPWR _00351_ sky130_fd_sc_hd__or2_1
X_09282_ _01360_ _01422_ VGND VGND VPWR VPWR _01423_ sky130_fd_sc_hd__and2_1
XFILLER_0_118_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07340__D _02149_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_142_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08233_ _00273_ _00276_ VGND VGND VPWR VPWR _00277_ sky130_fd_sc_hd__and2_1
XFILLER_0_62_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08164_ _04796_ _00207_ VGND VGND VPWR VPWR _00208_ sky130_fd_sc_hd__nor2_2
XFILLER_0_16_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07115_ _00563_ VGND VGND VPWR VPWR _00628_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__10402__A1 _05445_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08095_ _00138_ _02007_ _04928_ VGND VGND VPWR VPWR _00139_ sky130_fd_sc_hd__and3_1
XANTENNA__10402__B2 _05467_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_848 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_399 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_235 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_583 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08997_ _01107_ _01110_ VGND VGND VPWR VPWR _01111_ sky130_fd_sc_hd__or2b_1
X_07948_ _07037_ _07076_ VGND VGND VPWR VPWR _07077_ sky130_fd_sc_hd__and2_1
XANTENNA__10222__C _02029_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07879_ _06956_ _06959_ _07007_ VGND VGND VPWR VPWR _07008_ sky130_fd_sc_hd__a21o_1
XANTENNA__07334__A1 _02138_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08531__B1 _00379_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07334__B2 _00333_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09618_ _01582_ _01594_ VGND VGND VPWR VPWR _01791_ sky130_fd_sc_hd__nand2_1
X_10890_ _03182_ _03183_ VGND VGND VPWR VPWR _03185_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09549_ _01544_ _01554_ _01714_ VGND VGND VPWR VPWR _01715_ sky130_fd_sc_hd__a21o_1
XFILLER_0_66_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09087__B2 _01306_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12560_ _00390_ _04714_ _05020_ VGND VGND VPWR VPWR _05021_ sky130_fd_sc_hd__a21o_1
XFILLER_0_66_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11511_ _03849_ _03866_ VGND VGND VPWR VPWR _03867_ sky130_fd_sc_hd__nor2_1
XFILLER_0_80_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09739__B _01076_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12491_ _00613_ _03696_ _03729_ _00612_ VGND VGND VPWR VPWR _04945_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11350__A _03687_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14230_ _00206_ _00360_ VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__xor2_4
XFILLER_0_136_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11442_ _06964_ _02133_ _02459_ _00121_ VGND VGND VPWR VPWR _03791_ sky130_fd_sc_hd__a22o_1
XANTENNA__12394__A1 _00778_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12394__B2 _00782_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13591__B1 _02858_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14161_ _06752_ _06760_ VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__xnor2_4
X_11373_ _03713_ _03714_ VGND VGND VPWR VPWR _03715_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_22_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08062__A2 _06885_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10324_ _02561_ _02562_ VGND VGND VPWR VPWR _02563_ sky130_fd_sc_hd__and2b_1
X_13112_ _05624_ _05626_ _05627_ VGND VGND VPWR VPWR _05628_ sky130_fd_sc_hd__o21a_1
X_14092_ _05964_ _06685_ _06619_ _05959_ VGND VGND VPWR VPWR _06687_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_131_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13043_ _04579_ _04572_ VGND VGND VPWR VPWR _05552_ sky130_fd_sc_hd__or2b_1
X_10255_ _02485_ _02486_ _02483_ _02484_ VGND VGND VPWR VPWR _02488_ sky130_fd_sc_hd__o211a_1
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10186_ _02411_ VGND VGND VPWR VPWR _02413_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13945_ _06524_ _06525_ VGND VGND VPWR VPWR _06526_ sky130_fd_sc_hd__nand2_1
XANTENNA__07325__A1 _00464_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13876_ _06436_ _06445_ _06449_ VGND VGND VPWR VPWR _06451_ sky130_fd_sc_hd__and3_1
XFILLER_0_69_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12827_ _05312_ _05314_ VGND VGND VPWR VPWR _05315_ sky130_fd_sc_hd__nand2_1
XFILLER_0_146_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12758_ _00457_ _03738_ _04640_ _04639_ VGND VGND VPWR VPWR _05239_ sky130_fd_sc_hd__a31o_1
XFILLER_0_127_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11709_ _04054_ _04060_ VGND VGND VPWR VPWR _04085_ sky130_fd_sc_hd__nor2_1
XFILLER_0_126_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12689_ _04898_ _04909_ VGND VGND VPWR VPWR _05163_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12385__A1 _00778_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12385__B2 _00782_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07169__B net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09665__A _00843_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08920_ _00833_ _01025_ _01026_ VGND VGND VPWR VPWR _01027_ sky130_fd_sc_hd__and3_1
XFILLER_0_110_555 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07185__A _01208_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08851_ _03268_ net40 VGND VGND VPWR VPWR _00951_ sky130_fd_sc_hd__and2_1
X_07802_ _05170_ _05269_ _06930_ VGND VGND VPWR VPWR _06931_ sky130_fd_sc_hd__a21o_1
X_08782_ _00667_ _00704_ _00875_ VGND VGND VPWR VPWR _00876_ sky130_fd_sc_hd__o21ba_1
XANTENNA__07335__D _02971_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07733_ _06852_ _06861_ VGND VGND VPWR VPWR _06862_ sky130_fd_sc_hd__nand2_1
XANTENNA__08513__B1 _03938_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11435__A _03748_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07664_ _06494_ VGND VGND VPWR VPWR _06637_ sky130_fd_sc_hd__buf_4
XFILLER_0_67_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09403_ _01544_ _01554_ VGND VGND VPWR VPWR _01555_ sky130_fd_sc_hd__xor2_1
XFILLER_0_48_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07595_ _02029_ _05566_ _05753_ _05771_ VGND VGND VPWR VPWR _05879_ sky130_fd_sc_hd__a211o_1
XFILLER_0_62_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09334_ _01467_ _01478_ VGND VGND VPWR VPWR _01479_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09265_ _01067_ _01103_ _01102_ VGND VGND VPWR VPWR _01404_ sky130_fd_sc_hd__a21o_1
XFILLER_0_47_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08463__B _00526_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08216_ _00111_ _00116_ _00256_ _00259_ VGND VGND VPWR VPWR _00260_ sky130_fd_sc_hd__a211o_1
XFILLER_0_145_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09196_ _01326_ _01327_ VGND VGND VPWR VPWR _01329_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08147_ _06996_ _06995_ _06989_ VGND VGND VPWR VPWR _00191_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_114_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08078_ _06461_ _00121_ VGND VGND VPWR VPWR _00122_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13809__B _02189_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10514__A _02247_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07095__A _00399_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10040_ _01841_ _01844_ _02252_ VGND VGND VPWR VPWR _02253_ sky130_fd_sc_hd__o21a_1
XANTENNA__10233__B net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07823__A _00420_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11991_ _00530_ _01958_ _04393_ _03988_ VGND VGND VPWR VPWR _04395_ sky130_fd_sc_hd__a211o_1
XANTENNA__11345__A _03683_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07542__B _04939_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13730_ _06262_ _06287_ _06289_ VGND VGND VPWR VPWR _06290_ sky130_fd_sc_hd__o21a_1
X_10942_ _03221_ _03239_ _03240_ _03241_ VGND VGND VPWR VPWR _03242_ sky130_fd_sc_hd__a211o_1
XFILLER_0_86_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10311__B1 _00959_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13661_ _06016_ _06213_ VGND VGND VPWR VPWR _06214_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10873_ _03154_ _03164_ _03165_ VGND VGND VPWR VPWR _03166_ sky130_fd_sc_hd__o21a_1
XFILLER_0_128_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_840 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12612_ _05076_ _05077_ VGND VGND VPWR VPWR _05078_ sky130_fd_sc_hd__nand2_1
X_13592_ _06136_ _06137_ _01414_ _03785_ VGND VGND VPWR VPWR _06138_ sky130_fd_sc_hd__and4bb_1
XANTENNA__08654__A _00311_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_644 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12543_ _04998_ _04999_ _05001_ VGND VGND VPWR VPWR _05002_ sky130_fd_sc_hd__a21o_1
XFILLER_0_54_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12474_ _04913_ _04925_ VGND VGND VPWR VPWR _04926_ sky130_fd_sc_hd__xor2_2
XFILLER_0_123_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14213_ _01755_ _06801_ VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__nor2_4
XFILLER_0_62_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11425_ _03769_ _03771_ VGND VGND VPWR VPWR _03772_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08035__A2 _07075_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14144_ _06740_ _06741_ VGND VGND VPWR VPWR _06742_ sky130_fd_sc_hd__nor2_1
X_11356_ _03684_ VGND VGND VPWR VPWR _03697_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_104_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08820__C _00915_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10307_ _02355_ _02363_ _02544_ VGND VGND VPWR VPWR _02545_ sky130_fd_sc_hd__a21o_2
X_14075_ _06074_ _04013_ _06667_ VGND VGND VPWR VPWR _06668_ sky130_fd_sc_hd__and3_1
XTAP_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11287_ _03458_ _03467_ VGND VGND VPWR VPWR _03622_ sky130_fd_sc_hd__xor2_2
XANTENNA__10424__A net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13026_ _04573_ _05437_ VGND VGND VPWR VPWR _05534_ sky130_fd_sc_hd__nand2_1
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10238_ _02458_ _02469_ VGND VGND VPWR VPWR _02470_ sky130_fd_sc_hd__xnor2_2
XANTENNA__07546__A1 _02456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13735__A _00916_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10169_ _06965_ _00741_ _02014_ VGND VGND VPWR VPWR _02394_ sky130_fd_sc_hd__and3_1
XFILLER_0_83_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13454__B _02766_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xrebuffer19 _07039_ VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_107_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13928_ _06226_ _06228_ VGND VGND VPWR VPWR _06508_ sky130_fd_sc_hd__nor2_2
XFILLER_0_16_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13859_ _06401_ _06408_ VGND VGND VPWR VPWR _06432_ sky130_fd_sc_hd__xor2_1
XFILLER_0_9_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07380_ _03521_ VGND VGND VPWR VPWR _03532_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_146_227 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08283__B _02982_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09050_ _01042_ _01046_ VGND VGND VPWR VPWR _01169_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08001_ _00044_ VGND VGND VPWR VPWR _00045_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09223__A1 _00991_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_142_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09952_ net52 VGND VGND VPWR VPWR _02156_ sky130_fd_sc_hd__buf_2
XFILLER_0_0_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08903_ _00377_ _02993_ _00112_ _00268_ VGND VGND VPWR VPWR _01008_ sky130_fd_sc_hd__and4_1
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09883_ _02077_ _02079_ VGND VGND VPWR VPWR _02080_ sky130_fd_sc_hd__and2_1
XFILLER_0_110_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08834_ _00917_ _00744_ _00918_ _00931_ VGND VGND VPWR VPWR _00932_ sky130_fd_sc_hd__or4_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08765_ _00853_ _00856_ VGND VGND VPWR VPWR _00857_ sky130_fd_sc_hd__xor2_2
XFILLER_0_79_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07716_ _03598_ _06844_ VGND VGND VPWR VPWR _06845_ sky130_fd_sc_hd__and2_1
X_08696_ _00780_ VGND VGND VPWR VPWR _00782_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_68_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07647_ _06439_ VGND VGND VPWR VPWR _06450_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_94_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07578_ _05654_ _05665_ _05698_ VGND VGND VPWR VPWR _05709_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_82_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13811__C _01400_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12597__A1 _03740_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08905__C _06765_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09317_ _01337_ _01342_ _01460_ VGND VGND VPWR VPWR _01461_ sky130_fd_sc_hd__nor3_1
XANTENNA__12597__B2 _03707_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10509__A _02765_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09248_ _01384_ _01385_ VGND VGND VPWR VPWR _01386_ sky130_fd_sc_hd__or2_1
XFILLER_0_106_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09179_ _01115_ _01160_ VGND VGND VPWR VPWR _01310_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11210_ _02502_ _02541_ VGND VGND VPWR VPWR _03537_ sky130_fd_sc_hd__nor2_1
XFILLER_0_121_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12190_ _03608_ _03575_ _03610_ VGND VGND VPWR VPWR _04614_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_120_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__07776__A1 net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11141_ _03459_ _03460_ VGND VGND VPWR VPWR _03461_ sky130_fd_sc_hd__and2_2
XFILLER_0_9_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput66 net66 VGND VGND VPWR VPWR prod[10] sky130_fd_sc_hd__clkbuf_4
Xoutput77 net77 VGND VGND VPWR VPWR prod[20] sky130_fd_sc_hd__clkbuf_4
X_11072_ _03371_ _03383_ VGND VGND VPWR VPWR _03385_ sky130_fd_sc_hd__and2_1
Xoutput88 net88 VGND VGND VPWR VPWR prod[30] sky130_fd_sc_hd__clkbuf_4
Xoutput99 net99 VGND VGND VPWR VPWR prod[40] sky130_fd_sc_hd__clkbuf_4
X_10023_ _02210_ _02232_ VGND VGND VPWR VPWR _02234_ sky130_fd_sc_hd__nand2_1
XANTENNA__08649__A net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11974_ _04375_ _04373_ VGND VGND VPWR VPWR _04376_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09820__A1_N _03696_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13713_ _02427_ _02758_ _06264_ _05887_ _02726_ VGND VGND VPWR VPWR _06271_ sky130_fd_sc_hd__a32o_1
X_10925_ _03218_ _03222_ VGND VGND VPWR VPWR _03223_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_39_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13290__A _05810_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13644_ _06193_ _06194_ VGND VGND VPWR VPWR _06195_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08384__A _02467_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10856_ _06483_ _02857_ _03146_ VGND VGND VPWR VPWR _03148_ sky130_fd_sc_hd__and3_1
XFILLER_0_85_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13575_ _06009_ _05969_ _06018_ _05985_ VGND VGND VPWR VPWR _06119_ sky130_fd_sc_hd__and4_1
XFILLER_0_27_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10787_ _03063_ _03071_ VGND VGND VPWR VPWR _03072_ sky130_fd_sc_hd__and2b_1
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12526_ _04980_ _04981_ _04934_ VGND VGND VPWR VPWR _04984_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_54_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_444 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12457_ _04903_ _04904_ VGND VGND VPWR VPWR _04908_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_output91_A net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07728__A _00563_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11408_ _03749_ _03752_ _03753_ VGND VGND VPWR VPWR _03754_ sky130_fd_sc_hd__and3_1
X_12388_ _00784_ _00779_ _01586_ _01584_ VGND VGND VPWR VPWR _04832_ sky130_fd_sc_hd__nand4_1
XANTENNA__08964__B1 _00959_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14127_ _06722_ _06724_ VGND VGND VPWR VPWR _06725_ sky130_fd_sc_hd__nor2_1
XFILLER_0_22_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11339_ _02673_ VGND VGND VPWR VPWR _03678_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_120_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14058_ _06111_ VGND VGND VPWR VPWR _06650_ sky130_fd_sc_hd__inv_2
X_13009_ _04584_ _04575_ _04580_ VGND VGND VPWR VPWR _05515_ sky130_fd_sc_hd__or3_4
XANTENNA__09662__B _01741_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08559__A _00410_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08550_ _04312_ _00452_ _00451_ VGND VGND VPWR VPWR _00622_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_89_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07501_ _04851_ VGND VGND VPWR VPWR _04862_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_76_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08481_ _00527_ _00546_ VGND VGND VPWR VPWR _00547_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_134_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07432_ net42 VGND VGND VPWR VPWR _04103_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12579__A1 _00393_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10974__D _01400_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12579__B2 _00390_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07363_ _03257_ _03323_ VGND VGND VPWR VPWR _03345_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09102_ _01224_ _01225_ VGND VGND VPWR VPWR _01226_ sky130_fd_sc_hd__or2b_1
XANTENNA__07455__B1 _03004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07294_ _02521_ net152 VGND VGND VPWR VPWR _02587_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_72_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_504 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09033_ _01133_ _01148_ VGND VGND VPWR VPWR _01150_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_475 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_171 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09935_ _02127_ _00322_ net21 _02133_ VGND VGND VPWR VPWR _02137_ sky130_fd_sc_hd__and4_1
XFILLER_0_0_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09866_ _02012_ _02019_ VGND VGND VPWR VPWR _02062_ sky130_fd_sc_hd__nand2_1
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09380__B1 _01508_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08817_ _00742_ VGND VGND VPWR VPWR _00914_ sky130_fd_sc_hd__clkbuf_4
X_09797_ _03070_ _01585_ _01983_ _01986_ VGND VGND VPWR VPWR _01987_ sky130_fd_sc_hd__a22oi_1
XTAP_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08748_ _00664_ _00838_ VGND VGND VPWR VPWR _00839_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08679_ _00740_ _00762_ VGND VGND VPWR VPWR _00763_ sky130_fd_sc_hd__xnor2_4
XTAP_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12719__A _05193_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10710_ _02973_ _02984_ _02986_ VGND VGND VPWR VPWR _02987_ sky130_fd_sc_hd__a21oi_1
XTAP_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10293__A2 net49 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07694__B1 _06820_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11690_ _06819_ _00571_ net15 _06874_ VGND VGND VPWR VPWR _04064_ sky130_fd_sc_hd__a22oi_1
XTAP_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10641_ _02904_ _02906_ _02909_ VGND VGND VPWR VPWR _02911_ sky130_fd_sc_hd__nor3_1
XFILLER_0_64_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13360_ _05337_ _05352_ _05883_ VGND VGND VPWR VPWR _05884_ sky130_fd_sc_hd__a21oi_1
X_10572_ _02833_ _02834_ VGND VGND VPWR VPWR _02835_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_770 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12311_ _00607_ _00575_ _01664_ _00415_ VGND VGND VPWR VPWR _04747_ sky130_fd_sc_hd__a22o_1
X_13291_ _05712_ _05813_ VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__xor2_4
XFILLER_0_51_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12242_ _04665_ _04668_ _04670_ VGND VGND VPWR VPWR _04671_ sky130_fd_sc_hd__and3_1
XFILLER_0_121_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08370__C _00672_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12742__A1 _00779_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12742__B2 _00784_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12173_ _04555_ _04586_ _04594_ VGND VGND VPWR VPWR _04595_ sky130_fd_sc_hd__or3_4
XFILLER_0_48_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11124_ _03270_ _03297_ VGND VGND VPWR VPWR _03442_ sky130_fd_sc_hd__and2_1
X_11055_ _03296_ _03295_ VGND VGND VPWR VPWR _03366_ sky130_fd_sc_hd__or2b_1
XANTENNA__08379__A _02335_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09913__D _01254_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07283__A _02259_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10006_ _02213_ _02214_ VGND VGND VPWR VPWR _02216_ sky130_fd_sc_hd__and2_1
XANTENNA__09910__A2 _01955_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10421__B _02459_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10808__A1 _06494_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11957_ _06417_ _00138_ _02134_ _03681_ VGND VGND VPWR VPWR _04358_ sky130_fd_sc_hd__and4_1
XFILLER_0_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10908_ _03192_ _03199_ _03204_ VGND VGND VPWR VPWR _03205_ sky130_fd_sc_hd__or3_2
XFILLER_0_46_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11888_ _04271_ _04281_ VGND VGND VPWR VPWR _04282_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_39_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13627_ _06169_ _06173_ _06176_ VGND VGND VPWR VPWR _06177_ sky130_fd_sc_hd__a21oi_1
X_10839_ _03127_ _03128_ VGND VGND VPWR VPWR _03129_ sky130_fd_sc_hd__and2_1
XFILLER_0_109_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13558_ _06099_ _06100_ VGND VGND VPWR VPWR _06101_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12509_ _04962_ _04964_ VGND VGND VPWR VPWR _04965_ sky130_fd_sc_hd__and2b_1
XFILLER_0_140_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13489_ _06011_ _06013_ _01062_ _03699_ VGND VGND VPWR VPWR _06025_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_2_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12364__A _00741_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07981_ _00021_ _00024_ VGND VGND VPWR VPWR _00025_ sky130_fd_sc_hd__xor2_1
XFILLER_0_10_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09720_ _01900_ _01901_ VGND VGND VPWR VPWR _01902_ sky130_fd_sc_hd__nor2_1
XANTENNA__08289__A _00497_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09823__D net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07193__A _01120_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09651_ _01307_ _01625_ _01826_ VGND VGND VPWR VPWR _01827_ sky130_fd_sc_hd__a21o_2
XANTENNA__11427__B _06885_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07624__C _05742_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10331__B _04048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08602_ _00481_ _00470_ VGND VGND VPWR VPWR _00679_ sky130_fd_sc_hd__and2b_1
X_09582_ _01749_ _01750_ VGND VGND VPWR VPWR _01751_ sky130_fd_sc_hd__and2b_1
XFILLER_0_89_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08533_ _00601_ _00602_ VGND VGND VPWR VPWR _00603_ sky130_fd_sc_hd__or2_1
XANTENNA__11871__A1_N _00004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08468__A2 _06873_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13461__A2 _02722_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11443__A _06964_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08464_ _00508_ _00294_ _00336_ VGND VGND VPWR VPWR _00528_ sky130_fd_sc_hd__and3_1
XFILLER_0_37_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07415_ _03883_ _03905_ VGND VGND VPWR VPWR _03916_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08395_ _00441_ _00443_ _00450_ VGND VGND VPWR VPWR _00452_ sky130_fd_sc_hd__nand3_1
XFILLER_0_147_399 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07346_ _01044_ _00880_ net26 _03147_ VGND VGND VPWR VPWR _03158_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08752__A _00257_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07277_ _02357_ _02390_ VGND VGND VPWR VPWR _02401_ sky130_fd_sc_hd__and2_1
XFILLER_0_5_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09016_ _01129_ _01130_ VGND VGND VPWR VPWR _01132_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11527__A2 _01957_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12721__B _01108_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09918_ _02117_ VGND VGND VPWR VPWR _02119_ sky130_fd_sc_hd__clkbuf_4
X_09849_ _02041_ _02043_ VGND VGND VPWR VPWR _02044_ sky130_fd_sc_hd__xor2_4
X_12860_ _05273_ _05349_ VGND VGND VPWR VPWR _05351_ sky130_fd_sc_hd__nand2_1
XTAP_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11811_ _06428_ _03748_ _04196_ VGND VGND VPWR VPWR _04197_ sky130_fd_sc_hd__and3_1
XTAP_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12791_ _05273_ _05274_ VGND VGND VPWR VPWR _05275_ sky130_fd_sc_hd__or2_1
XTAP_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11353__A _02246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11742_ _04117_ _04119_ _04120_ VGND VGND VPWR VPWR _04121_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11673_ _06733_ _03938_ _04042_ _04043_ VGND VGND VPWR VPWR _04045_ sky130_fd_sc_hd__o2bb2a_1
XTAP_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13412_ _05937_ _05940_ VGND VGND VPWR VPWR _05941_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_36_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10018__A2 _00376_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10624_ _02881_ _02890_ _02891_ VGND VGND VPWR VPWR _02892_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_52_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08662__A _00157_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13343_ _05854_ _05336_ _05864_ VGND VGND VPWR VPWR _05865_ sky130_fd_sc_hd__and3_1
XFILLER_0_122_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10555_ _02814_ _02815_ _00095_ _01933_ VGND VGND VPWR VPWR _02816_ sky130_fd_sc_hd__and4b_1
XFILLER_0_134_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13274_ _05784_ _05793_ _05797_ VGND VGND VPWR VPWR _05798_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_59_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10486_ _02734_ _02738_ _02739_ VGND VGND VPWR VPWR _02741_ sky130_fd_sc_hd__and3_1
XFILLER_0_32_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12225_ _00375_ _03744_ _04650_ _04651_ VGND VGND VPWR VPWR _04652_ sky130_fd_sc_hd__a31o_1
XANTENNA__09493__A _01372_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09592__B1 net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12156_ _02699_ VGND VGND VPWR VPWR _04577_ sky130_fd_sc_hd__inv_2
XFILLER_0_102_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11107_ _02562_ _02577_ VGND VGND VPWR VPWR _03424_ sky130_fd_sc_hd__and2_1
X_12087_ _04346_ _04351_ _04421_ VGND VGND VPWR VPWR _04501_ sky130_fd_sc_hd__o21a_1
X_11038_ net7 _00373_ VGND VGND VPWR VPWR _03348_ sky130_fd_sc_hd__nand2_1
XANTENNA__08259__D _04928_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13462__B _02735_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12989_ _05431_ _03611_ VGND VGND VPWR VPWR _05493_ sky130_fd_sc_hd__xnor2_4
XANTENNA__12359__A _00742_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13443__A2 _02766_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07200_ _01328_ _01547_ VGND VGND VPWR VPWR _01558_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08180_ _00216_ _00223_ VGND VGND VPWR VPWR _00224_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_55_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07131_ _00781_ _00792_ VGND VGND VPWR VPWR _00803_ sky130_fd_sc_hd__xnor2_2
XANTENNA__11710__B _00915_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10607__A _00158_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_507 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07188__A _01350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07594__C1 _05566_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11438__A _00843_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07964_ _07009_ _07015_ VGND VGND VPWR VPWR _00008_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12260__C _01180_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09703_ _01709_ _01882_ VGND VGND VPWR VPWR _01883_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07895_ _07022_ _07023_ VGND VGND VPWR VPWR _07024_ sky130_fd_sc_hd__nor2_1
X_09634_ _01197_ _04510_ net18 VGND VGND VPWR VPWR _01808_ sky130_fd_sc_hd__and3_1
XANTENNA__07651__A _06483_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09565_ _01726_ _01727_ _01729_ _01730_ VGND VGND VPWR VPWR _01732_ sky130_fd_sc_hd__o22a_1
XFILLER_0_78_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08516_ _00581_ _00582_ _00422_ _00425_ VGND VGND VPWR VPWR _00585_ sky130_fd_sc_hd__a211oi_1
X_09496_ _01284_ net49 _01548_ _01655_ VGND VGND VPWR VPWR _01657_ sky130_fd_sc_hd__a31o_1
XFILLER_0_37_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08447_ _00309_ _00313_ _00507_ VGND VGND VPWR VPWR _00510_ sky130_fd_sc_hd__nor3_1
XFILLER_0_136_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11901__A _02280_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08378_ _00432_ _00433_ VGND VGND VPWR VPWR _00434_ sky130_fd_sc_hd__nor2_1
XFILLER_0_135_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07329_ _02960_ VGND VGND VPWR VPWR _02971_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_33_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07098__A _00431_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10340_ _02233_ _02376_ _02580_ VGND VGND VPWR VPWR _02581_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_21_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10271_ _02303_ _02308_ VGND VGND VPWR VPWR _02505_ sky130_fd_sc_hd__nand2_1
X_12010_ _04337_ _04415_ VGND VGND VPWR VPWR _04416_ sky130_fd_sc_hd__and2_1
XANTENNA__07826__A _01076_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07545__B _00399_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13961_ _06543_ VGND VGND VPWR VPWR _06544_ sky130_fd_sc_hd__inv_2
X_12912_ _05406_ _05407_ VGND VGND VPWR VPWR _05408_ sky130_fd_sc_hd__nor2_1
X_13892_ _06456_ _06460_ _06467_ _06459_ VGND VGND VPWR VPWR _06468_ sky130_fd_sc_hd__o22a_1
X_12843_ _05326_ _05331_ VGND VGND VPWR VPWR _05332_ sky130_fd_sc_hd__xor2_1
XTAP_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_620 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12633__B1 _02723_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12774_ _05254_ _05255_ VGND VGND VPWR VPWR _05256_ sky130_fd_sc_hd__or2b_1
XTAP_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08095__C _04928_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11725_ _04083_ _04101_ VGND VGND VPWR VPWR _04102_ sky130_fd_sc_hd__nor2_1
XFILLER_0_138_163 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11811__A _06428_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11656_ _04011_ _03859_ _04009_ VGND VGND VPWR VPWR _04027_ sky130_fd_sc_hd__or3_1
XFILLER_0_36_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11739__A2 _01188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10607_ _00158_ _01059_ VGND VGND VPWR VPWR _02874_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11587_ _03943_ _03947_ _03950_ VGND VGND VPWR VPWR _03951_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13326_ _05647_ _05663_ _05829_ _05846_ VGND VGND VPWR VPWR _05848_ sky130_fd_sc_hd__a31o_1
XFILLER_0_122_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07812__B1 _06820_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10538_ _00293_ _02725_ _02728_ _03015_ VGND VGND VPWR VPWR _02798_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13257_ _05758_ _05781_ VGND VGND VPWR VPWR _05782_ sky130_fd_sc_hd__and2_1
X_10469_ _02721_ VGND VGND VPWR VPWR _02722_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_86_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09935__B _00322_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07736__A _00420_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12208_ _01518_ _01954_ _02135_ _00375_ VGND VGND VPWR VPWR _04634_ sky130_fd_sc_hd__a22oi_1
XANTENNA__10175__A1 _00101_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13188_ _05696_ _05711_ VGND VGND VPWR VPWR _05712_ sky130_fd_sc_hd__xnor2_4
XANTENNA__10175__B2 net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12139_ _02596_ _02644_ VGND VGND VPWR VPWR _04558_ sky130_fd_sc_hd__nor2_1
XANTENNA__09868__A1 _06873_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09868__B2 _06875_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10478__A2 _02726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07680_ net1 net35 net34 net12 VGND VGND VPWR VPWR _06797_ sky130_fd_sc_hd__a22o_1
XANTENNA__08540__A1 _04268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08286__B _00094_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09350_ _01495_ _01496_ VGND VGND VPWR VPWR _01497_ sky130_fd_sc_hd__xor2_1
XFILLER_0_87_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08301_ _04004_ _00349_ VGND VGND VPWR VPWR _00350_ sky130_fd_sc_hd__xnor2_4
X_09281_ _01365_ _01421_ VGND VGND VPWR VPWR _01422_ sky130_fd_sc_hd__xor2_1
XFILLER_0_142_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09398__A _01372_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08232_ _00274_ _00275_ VGND VGND VPWR VPWR _00276_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_62_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08163_ _04774_ _04785_ VGND VGND VPWR VPWR _00207_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07114_ _00552_ _00606_ VGND VGND VPWR VPWR _00617_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_113_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10402__A2 _01177_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08094_ _05478_ VGND VGND VPWR VPWR _00138_ sky130_fd_sc_hd__buf_2
XFILLER_0_101_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07646__A _05478_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_595 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08996_ _00464_ _01108_ _01106_ VGND VGND VPWR VPWR _01110_ sky130_fd_sc_hd__a21o_1
X_07947_ net165 _07075_ VGND VGND VPWR VPWR _07076_ sky130_fd_sc_hd__xor2_1
X_07878_ _01230_ _06744_ _06957_ VGND VGND VPWR VPWR _07007_ sky130_fd_sc_hd__and3_1
XANTENNA__08477__A _07004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08531__A1 _02259_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07334__A2 _00410_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07381__A _03532_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08531__B2 _02171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09617_ _01787_ _01789_ VGND VGND VPWR VPWR _01790_ sky130_fd_sc_hd__nand2_1
X_09548_ _01544_ _01554_ _01500_ VGND VGND VPWR VPWR _01714_ sky130_fd_sc_hd__o21a_1
XANTENNA__09087__A2 _00730_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09479_ _01432_ _01638_ VGND VGND VPWR VPWR _01639_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11510_ _03846_ _03848_ VGND VGND VPWR VPWR _03866_ sky130_fd_sc_hd__and2_1
XFILLER_0_81_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12490_ _04941_ _04943_ VGND VGND VPWR VPWR _04944_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_80_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11441_ _03754_ _03787_ _03752_ VGND VGND VPWR VPWR _03790_ sky130_fd_sc_hd__a21bo_1
Xwire136 _06487_ VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__buf_1
XFILLER_0_18_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_142 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12394__A2 _00413_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14160_ _06756_ _06757_ _06758_ _06759_ _06643_ VGND VGND VPWR VPWR _06760_ sky130_fd_sc_hd__a311oi_4
XANTENNA__13591__A1 _01250_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11372_ _01155_ _03697_ VGND VGND VPWR VPWR _03714_ sky130_fd_sc_hd__nand2_2
XFILLER_0_61_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13591__B2 _01181_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13111_ _05605_ _05623_ VGND VGND VPWR VPWR _05627_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10323_ _02214_ _02546_ _02547_ _02560_ VGND VGND VPWR VPWR _02562_ sky130_fd_sc_hd__a31o_1
XFILLER_0_131_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_575 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14091_ _05961_ _06685_ VGND VGND VPWR VPWR _06686_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13042_ _05550_ _04605_ _02589_ VGND VGND VPWR VPWR _05551_ sky130_fd_sc_hd__mux2_1
X_10254_ _02483_ _02484_ _02485_ _02486_ VGND VGND VPWR VPWR _02487_ sky130_fd_sc_hd__a211oi_2
XANTENNA__11354__B1 _03690_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10185_ _06821_ net13 _00730_ _03499_ VGND VGND VPWR VPWR _02411_ sky130_fd_sc_hd__a22o_1
XANTENNA__09771__A _01957_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13944_ _06453_ _06478_ VGND VGND VPWR VPWR _06525_ sky130_fd_sc_hd__xor2_2
XANTENNA__07325__A2 _00530_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13875_ _06447_ _06448_ VGND VGND VPWR VPWR _06449_ sky130_fd_sc_hd__or2_1
XFILLER_0_88_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12826_ _05311_ _05140_ _05218_ VGND VGND VPWR VPWR _05314_ sky130_fd_sc_hd__nand3_1
XFILLER_0_96_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12757_ _05235_ _05237_ VGND VGND VPWR VPWR _05238_ sky130_fd_sc_hd__xor2_1
XTAP_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11708_ _04041_ _04046_ _04053_ VGND VGND VPWR VPWR _04084_ sky130_fd_sc_hd__and3_1
XFILLER_0_127_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12688_ _04926_ _05033_ _05034_ VGND VGND VPWR VPWR _05162_ sky130_fd_sc_hd__a21o_1
XFILLER_0_127_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11260__B _03527_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09011__A _00003_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11639_ _03875_ _04006_ _04007_ VGND VGND VPWR VPWR _04008_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_142_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12385__A2 _00571_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07169__C _01197_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13309_ _05814_ _05826_ VGND VGND VPWR VPWR _05831_ sky130_fd_sc_hd__and2_1
XANTENNA__09665__B _00670_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12372__A _00914_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08850_ _02664_ net40 _00768_ _00767_ VGND VGND VPWR VPWR _00950_ sky130_fd_sc_hd__a31o_1
X_07801_ _05170_ _05269_ _05082_ VGND VGND VPWR VPWR _06930_ sky130_fd_sc_hd__o21ba_1
X_08781_ _00667_ _00704_ _00666_ VGND VGND VPWR VPWR _00875_ sky130_fd_sc_hd__a21boi_1
X_07732_ _06859_ _06860_ VGND VGND VPWR VPWR _06861_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08513__A1 _01295_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08513__B2 _01405_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07663_ _06428_ VGND VGND VPWR VPWR _06626_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_95_808 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09402_ _01552_ _01553_ VGND VGND VPWR VPWR _01554_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07594_ _05753_ _05771_ _02029_ _05566_ VGND VGND VPWR VPWR _05868_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_62_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09333_ _01476_ _01477_ VGND VGND VPWR VPWR _01478_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11451__A _06964_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09264_ _01398_ _01402_ VGND VGND VPWR VPWR _01403_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_118_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09559__C _00654_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08215_ _01383_ _01350_ _00257_ _00258_ VGND VGND VPWR VPWR _00259_ sky130_fd_sc_hd__and4_1
XFILLER_0_118_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09195_ _01325_ _01324_ VGND VGND VPWR VPWR _01327_ sky130_fd_sc_hd__and2b_1
XFILLER_0_62_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_199 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08146_ _06989_ _06996_ _06995_ VGND VGND VPWR VPWR _00190_ sky130_fd_sc_hd__or3_4
XFILLER_0_31_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13378__A _01664_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08077_ _06874_ VGND VGND VPWR VPWR _00121_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__13809__C _01954_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10514__B _02765_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10233__C _00322_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09591__A _06818_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08979_ _03268_ _04026_ VGND VGND VPWR VPWR _01091_ sky130_fd_sc_hd__nand2_1
XANTENNA__07823__B net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11990_ _04393_ _03988_ _00530_ _01958_ VGND VGND VPWR VPWR _04394_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_98_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10941_ _03215_ _03219_ _03207_ VGND VGND VPWR VPWR _03241_ sky130_fd_sc_hd__o21a_1
XANTENNA__10311__A1 _02971_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08000__A _03059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10311__B2 _00366_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13660_ _01415_ _01958_ _06078_ _01108_ VGND VGND VPWR VPWR _06213_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_39_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10872_ _03145_ _03148_ VGND VGND VPWR VPWR _03165_ sky130_fd_sc_hd__xor2_1
XFILLER_0_38_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12611_ _00389_ _00393_ _01060_ _01412_ VGND VGND VPWR VPWR _05077_ sky130_fd_sc_hd__and4_1
XFILLER_0_94_852 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13591_ _01250_ _02856_ _02858_ _01181_ VGND VGND VPWR VPWR _06137_ sky130_fd_sc_hd__a22oi_1
XANTENNA__08654__B _00734_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11361__A _00843_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12542_ _04998_ _04999_ _05000_ VGND VGND VPWR VPWR _05001_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_109_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12473_ _04921_ _04923_ _04924_ VGND VGND VPWR VPWR _04925_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_108_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14212_ _00464_ _02138_ _00344_ _02051_ VGND VGND VPWR VPWR _06801_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_22_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11424_ _03747_ _03770_ VGND VGND VPWR VPWR _03771_ sky130_fd_sc_hd__and2_1
XANTENNA__09766__A net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14143_ _06739_ _06736_ VGND VGND VPWR VPWR _06741_ sky130_fd_sc_hd__and2b_1
X_11355_ _03693_ _03694_ _01312_ _03684_ VGND VGND VPWR VPWR _03695_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_1_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10306_ _02355_ _02363_ _02374_ VGND VGND VPWR VPWR _02544_ sky130_fd_sc_hd__o21ba_1
X_14074_ _06075_ _06077_ _06078_ _02743_ _06107_ VGND VGND VPWR VPWR _06667_ sky130_fd_sc_hd__a41o_1
XFILLER_0_131_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08820__D _00916_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11286_ _03619_ _03615_ VGND VGND VPWR VPWR _03621_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13025_ _05516_ _05531_ VGND VGND VPWR VPWR _05532_ sky130_fd_sc_hd__or2b_2
X_10237_ _02466_ _02468_ VGND VGND VPWR VPWR _02469_ sky130_fd_sc_hd__nand2_1
XANTENNA__07546__A2 _00399_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10168_ _02063_ _02064_ _02065_ VGND VGND VPWR VPWR _02393_ sky130_fd_sc_hd__and3_1
XANTENNA__13735__B _02730_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11536__A _06819_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10099_ _02315_ _02316_ VGND VGND VPWR VPWR _02317_ sky130_fd_sc_hd__xor2_1
X_13927_ net134 _06506_ VGND VGND VPWR VPWR _06507_ sky130_fd_sc_hd__or2_2
XFILLER_0_16_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13858_ _06423_ _06430_ VGND VGND VPWR VPWR _06431_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_707 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08845__A _00563_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12809_ _05275_ _05294_ VGND VGND VPWR VPWR _05295_ sky130_fd_sc_hd__xor2_1
X_13789_ _06343_ _06353_ _06354_ VGND VGND VPWR VPWR _06355_ sky130_fd_sc_hd__a21o_1
XFILLER_0_146_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08283__C _06873_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08000_ _03059_ _02040_ _04917_ _04939_ VGND VGND VPWR VPWR _00044_ sky130_fd_sc_hd__and4_1
XFILLER_0_13_602 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_810 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07196__A _00420_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09951_ _01339_ _01410_ _01924_ _01923_ VGND VGND VPWR VPWR _02155_ sky130_fd_sc_hd__a31o_1
XFILLER_0_111_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07627__C _01996_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08902_ _01005_ _01006_ VGND VGND VPWR VPWR _01007_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09882_ _02078_ VGND VGND VPWR VPWR _02079_ sky130_fd_sc_hd__inv_2
XANTENNA__11869__A1 _06775_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11869__B2 _00575_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08833_ _00929_ _00930_ VGND VGND VPWR VPWR _00931_ sky130_fd_sc_hd__nor2_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08764_ _00469_ _00492_ _00854_ _00855_ VGND VGND VPWR VPWR _00856_ sky130_fd_sc_hd__a31o_1
X_07715_ _06842_ _06843_ VGND VGND VPWR VPWR _06844_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12294__A1 _03414_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08695_ _04180_ VGND VGND VPWR VPWR _00780_ sky130_fd_sc_hd__buf_2
XFILLER_0_73_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07646_ _05478_ VGND VGND VPWR VPWR _06439_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08755__A _06637_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07577_ _05676_ _05687_ VGND VGND VPWR VPWR _05698_ sky130_fd_sc_hd__and2_1
XANTENNA__13811__D _03683_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09316_ _01457_ _01458_ VGND VGND VPWR VPWR _01460_ sky130_fd_sc_hd__xor2_1
XANTENNA__12597__A2 _01411_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10188__A1_N _00486_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08905__D _00095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09247_ _02664_ _02719_ _00780_ _00777_ VGND VGND VPWR VPWR _01385_ sky130_fd_sc_hd__and4_2
XFILLER_0_118_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__08670__B1 _03718_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09178_ _01307_ _01308_ VGND VGND VPWR VPWR _01309_ sky130_fd_sc_hd__nor2_4
XFILLER_0_90_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08129_ _00075_ _00076_ VGND VGND VPWR VPWR _00173_ sky130_fd_sc_hd__nor2_1
XANTENNA__07776__A2 net6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11140_ _03305_ _03447_ VGND VGND VPWR VPWR _03460_ sky130_fd_sc_hd__xor2_2
XANTENNA__10780__A1 _06637_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput67 net67 VGND VGND VPWR VPWR prod[11] sky130_fd_sc_hd__clkbuf_4
Xoutput78 net78 VGND VGND VPWR VPWR prod[21] sky130_fd_sc_hd__buf_2
X_11071_ _03371_ _03383_ VGND VGND VPWR VPWR _03384_ sky130_fd_sc_hd__nor2_1
Xoutput89 net89 VGND VGND VPWR VPWR prod[31] sky130_fd_sc_hd__buf_2
X_10022_ _02210_ _02232_ VGND VGND VPWR VPWR _02233_ sky130_fd_sc_hd__or2_4
XFILLER_0_98_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11973_ _04308_ _04310_ VGND VGND VPWR VPWR _04375_ sky130_fd_sc_hd__and2_1
XFILLER_0_86_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10924_ _03215_ _03216_ VGND VGND VPWR VPWR _03222_ sky130_fd_sc_hd__or2_1
X_13712_ _06256_ _06269_ VGND VGND VPWR VPWR _06270_ sky130_fd_sc_hd__or2_1
XFILLER_0_85_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13643_ _06133_ _06167_ VGND VGND VPWR VPWR _06194_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_39_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10855_ _06461_ _02855_ VGND VGND VPWR VPWR _03146_ sky130_fd_sc_hd__nand2_1
XANTENNA__08384__B _00381_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13574_ _05992_ _06117_ VGND VGND VPWR VPWR _06118_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10786_ _03068_ _03069_ VGND VGND VPWR VPWR _03071_ sky130_fd_sc_hd__and2_1
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11796__B1 _02673_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12525_ _04934_ _04980_ _04981_ VGND VGND VPWR VPWR _04982_ sky130_fd_sc_hd__or3_1
XFILLER_0_82_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12456_ _04765_ _04766_ VGND VGND VPWR VPWR _04907_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_124_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11548__B1 _02120_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11407_ _00257_ _03750_ _03748_ _00670_ VGND VGND VPWR VPWR _03753_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07728__B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_49 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12387_ _00374_ _01584_ _04828_ _04830_ VGND VGND VPWR VPWR _04831_ sky130_fd_sc_hd__a31o_1
XFILLER_0_1_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14126_ _06720_ _06721_ VGND VGND VPWR VPWR _06724_ sky130_fd_sc_hd__and2_1
XANTENNA__08964__A1 _01076_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output84_A net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08964__B2 _03587_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11338_ _02793_ _03675_ _03676_ VGND VGND VPWR VPWR _03677_ sky130_fd_sc_hd__or3b_1
XFILLER_0_120_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14057_ _06238_ _06609_ VGND VGND VPWR VPWR _06649_ sky130_fd_sc_hd__or2_2
X_11269_ _03597_ _03601_ VGND VGND VPWR VPWR _03602_ sky130_fd_sc_hd__xor2_2
XFILLER_0_120_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13008_ _03578_ _04602_ _04606_ VGND VGND VPWR VPWR _05514_ sky130_fd_sc_hd__nand3_1
XANTENNA__07744__A _06819_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08559__B _00544_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13481__A _01062_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07500_ net5 VGND VGND VPWR VPWR _04851_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__09000__B1_N _01032_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08480_ _00542_ _00545_ VGND VGND VPWR VPWR _00546_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07431_ _04081_ _04048_ VGND VGND VPWR VPWR _04092_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12579__A2 _02758_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07362_ _03257_ _03323_ VGND VGND VPWR VPWR _03334_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09101_ _00932_ _01223_ _01190_ VGND VGND VPWR VPWR _01225_ sky130_fd_sc_hd__nand3_1
XFILLER_0_17_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07455__A1 _02018_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_143_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07293_ _02554_ _02565_ VGND VGND VPWR VPWR _02576_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07455__B2 _02040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09032_ _01133_ _01148_ VGND VGND VPWR VPWR _01149_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_763 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10064__B _02278_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09934_ _02138_ _01954_ _02135_ _00333_ VGND VGND VPWR VPWR _02136_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09865_ _06765_ _06775_ _03707_ _03740_ VGND VGND VPWR VPWR _02060_ sky130_fd_sc_hd__nand4_2
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09380__B2 _02116_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08816_ _00910_ _00911_ VGND VGND VPWR VPWR _00913_ sky130_fd_sc_hd__or2_2
XFILLER_0_99_229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09796_ _01984_ VGND VGND VPWR VPWR _01986_ sky130_fd_sc_hd__inv_2
XANTENNA__07930__A2 net6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08747_ _00806_ _00837_ VGND VGND VPWR VPWR _00838_ sky130_fd_sc_hd__xnor2_1
XTAP_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13391__A _01518_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08678_ _00751_ _00761_ VGND VGND VPWR VPWR _00762_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_68_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07694__A1 _01076_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07629_ _06230_ _06241_ VGND VGND VPWR VPWR _06252_ sky130_fd_sc_hd__nor2_1
XTAP_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07694__B2 _01120_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10640_ _02904_ _02906_ _02909_ VGND VGND VPWR VPWR _02910_ sky130_fd_sc_hd__o21a_1
XFILLER_0_119_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07446__A1 _01284_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10571_ _00399_ _03015_ _01934_ _02169_ VGND VGND VPWR VPWR _02834_ sky130_fd_sc_hd__and4_1
XFILLER_0_146_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08932__B _01039_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12310_ _04733_ _04745_ VGND VGND VPWR VPWR _04746_ sky130_fd_sc_hd__nor2_1
XANTENNA__07829__A _01120_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13290_ _05810_ _05811_ _05812_ VGND VGND VPWR VPWR _05813_ sky130_fd_sc_hd__nand3_2
XFILLER_0_51_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12241_ _04656_ _04669_ VGND VGND VPWR VPWR _04670_ sky130_fd_sc_hd__nor2_1
XFILLER_0_121_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08370__D net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12742__A2 _01953_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12172_ _04591_ _04552_ _04593_ VGND VGND VPWR VPWR _04594_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10753__A1 _00399_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11123_ _03419_ _03438_ _03439_ _03440_ VGND VGND VPWR VPWR _03441_ sky130_fd_sc_hd__a211o_1
XFILLER_0_101_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11054_ _03335_ _03364_ VGND VGND VPWR VPWR _03365_ sky130_fd_sc_hd__and2_1
XANTENNA__08379__B _00389_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10005_ _05203_ _04598_ _00782_ _00613_ VGND VGND VPWR VPWR _02214_ sky130_fd_sc_hd__nand4_1
XFILLER_0_64_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output122_A net122 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10808__A2 _01934_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11956_ _04353_ _04354_ _04355_ VGND VGND VPWR VPWR _04357_ sky130_fd_sc_hd__nand3_2
XFILLER_0_86_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10907_ _03201_ _03203_ VGND VGND VPWR VPWR _03204_ sky130_fd_sc_hd__nor2_1
X_11887_ _04278_ _04280_ VGND VGND VPWR VPWR _04281_ sky130_fd_sc_hd__or2b_1
XFILLER_0_67_660 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13626_ _06048_ _06174_ VGND VGND VPWR VPWR _06176_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10838_ _03119_ _03122_ VGND VGND VPWR VPWR _03128_ sky130_fd_sc_hd__xor2_1
XFILLER_0_55_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13557_ _06091_ _06097_ VGND VGND VPWR VPWR _06100_ sky130_fd_sc_hd__or2_1
XFILLER_0_70_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10769_ _02935_ _03001_ _03051_ VGND VGND VPWR VPWR _03052_ sky130_fd_sc_hd__o21bai_4
XFILLER_0_89_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07739__A _01284_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12508_ _04957_ _04963_ VGND VGND VPWR VPWR _04964_ sky130_fd_sc_hd__xnor2_1
X_13488_ _06022_ _06023_ VGND VGND VPWR VPWR _06024_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_81_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12364__B _00457_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12439_ _04767_ _04768_ VGND VGND VPWR VPWR _04888_ sky130_fd_sc_hd__or2_1
XFILLER_0_112_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14109_ _06703_ _06704_ VGND VGND VPWR VPWR _06705_ sky130_fd_sc_hd__nor2_1
XANTENNA__13476__A _01414_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07980_ _00022_ _00023_ VGND VGND VPWR VPWR _00024_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08289__B _00151_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07193__B _01470_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09650_ _01563_ _01623_ VGND VGND VPWR VPWR _01826_ sky130_fd_sc_hd__and2_1
XANTENNA__11427__C _01180_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07624__D _02664_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08601_ _00676_ _00677_ VGND VGND VPWR VPWR _00678_ sky130_fd_sc_hd__or2_1
X_09581_ _01465_ _01723_ _01748_ VGND VGND VPWR VPWR _01750_ sky130_fd_sc_hd__nand3_1
XFILLER_0_145_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08532_ _02105_ _02149_ _04037_ _04048_ VGND VGND VPWR VPWR _00602_ sky130_fd_sc_hd__and4_1
XFILLER_0_89_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07125__B1 net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08463_ _00519_ _00526_ VGND VGND VPWR VPWR _00527_ sky130_fd_sc_hd__nand2_1
XANTENNA__11443__B _00121_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07414_ _02127_ _03894_ VGND VGND VPWR VPWR _03905_ sky130_fd_sc_hd__nand2_1
X_08394_ _00441_ _00443_ _00450_ VGND VGND VPWR VPWR _00451_ sky130_fd_sc_hd__a21o_1
XFILLER_0_70_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07345_ net61 VGND VGND VPWR VPWR _03147_ sky130_fd_sc_hd__buf_2
XFILLER_0_128_592 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07649__A _06461_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07276_ _02379_ VGND VGND VPWR VPWR _02390_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_242 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09015_ _01119_ _01121_ _01128_ VGND VGND VPWR VPWR _01130_ sky130_fd_sc_hd__or3_1
XFILLER_0_115_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_584 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07384__A _00431_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09917_ _01361_ _02117_ _01960_ _00159_ VGND VGND VPWR VPWR _02118_ sky130_fd_sc_hd__a22o_1
X_09848_ _01760_ _02042_ VGND VGND VPWR VPWR _02043_ sky130_fd_sc_hd__or2b_2
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09779_ _01197_ _04510_ _01246_ net19 VGND VGND VPWR VPWR _01967_ sky130_fd_sc_hd__and4_1
XTAP_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ _06439_ _03750_ VGND VGND VPWR VPWR _04196_ sky130_fd_sc_hd__nand2_1
XTAP_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12790_ _05097_ _05272_ VGND VGND VPWR VPWR _05274_ sky130_fd_sc_hd__and2_1
XTAP_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11353__B _02249_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11741_ _04113_ _04116_ VGND VGND VPWR VPWR _04120_ sky130_fd_sc_hd__nand2_1
XTAP_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10671__B1 _02304_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11672_ _04042_ _04043_ _06733_ net11 VGND VGND VPWR VPWR _04044_ sky130_fd_sc_hd__and4bb_1
XTAP_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_855 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13411_ _05938_ _05939_ VGND VGND VPWR VPWR _05940_ sky130_fd_sc_hd__nand2_1
X_10623_ _02880_ _02878_ VGND VGND VPWR VPWR _02891_ sky130_fd_sc_hd__and2b_1
XFILLER_0_107_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08662__B _00741_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07559__A _05456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13342_ _05861_ _05863_ VGND VGND VPWR VPWR _05864_ sky130_fd_sc_hd__or2_1
X_10554_ _02993_ _02168_ _02723_ _00377_ VGND VGND VPWR VPWR _02815_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13273_ _05600_ _05506_ _05796_ VGND VGND VPWR VPWR _05797_ sky130_fd_sc_hd__a21oi_1
X_10485_ _02247_ _02736_ _02737_ _01473_ VGND VGND VPWR VPWR _02739_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09774__A _00322_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12224_ _00783_ _00778_ _01248_ _02117_ VGND VGND VPWR VPWR _04651_ sky130_fd_sc_hd__and4_1
XANTENNA__09592__A1 _06818_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12155_ _04567_ _04573_ _04574_ VGND VGND VPWR VPWR _04575_ sky130_fd_sc_hd__a21oi_4
XANTENNA__09493__B net50 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09592__B2 _06820_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11106_ _07040_ _01066_ VGND VGND VPWR VPWR _03423_ sky130_fd_sc_hd__and2_1
X_12086_ _04497_ _04498_ VGND VGND VPWR VPWR _04500_ sky130_fd_sc_hd__nor2_2
X_11037_ _03337_ _03336_ VGND VGND VPWR VPWR _03347_ sky130_fd_sc_hd__and2b_1
XFILLER_0_91_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12988_ _05472_ _05491_ VGND VGND VPWR VPWR _05492_ sky130_fd_sc_hd__and2_1
XANTENNA__12359__B _00605_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11939_ _04258_ _04260_ _04336_ VGND VGND VPWR VPWR _04338_ sky130_fd_sc_hd__nor3_1
XFILLER_0_24_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13609_ _05951_ _06156_ VGND VGND VPWR VPWR _06157_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07130_ net30 net33 VGND VGND VPWR VPWR _00792_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07469__A _00573_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10607__B _01059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07188__B _01361_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_390 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11719__A _00262_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07594__B1 _02029_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11438__B _03783_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07963_ _00005_ _00006_ VGND VGND VPWR VPWR _00007_ sky130_fd_sc_hd__nor2_1
XANTENNA__10342__B _02582_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09702_ _01880_ _01881_ VGND VGND VPWR VPWR _01882_ sky130_fd_sc_hd__or2b_1
XANTENNA__12260__D _01249_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07894_ net28 net29 _06818_ net34 VGND VGND VPWR VPWR _07023_ sky130_fd_sc_hd__and4_1
XANTENNA__07346__B1 net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09633_ _01773_ _01806_ VGND VGND VPWR VPWR _01807_ sky130_fd_sc_hd__xnor2_2
XANTENNA__13419__B1 _01252_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09564_ _01726_ _01727_ _01729_ _01730_ VGND VGND VPWR VPWR _01731_ sky130_fd_sc_hd__nor4_1
XANTENNA__11792__A2_N net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08515_ _00422_ _00425_ _00581_ _00582_ VGND VGND VPWR VPWR _00583_ sky130_fd_sc_hd__o211a_1
X_09495_ _00431_ _04169_ net50 net51 VGND VGND VPWR VPWR _01655_ sky130_fd_sc_hd__and4_1
XFILLER_0_93_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08446_ _00309_ net145 _00507_ VGND VGND VPWR VPWR _00509_ sky130_fd_sc_hd__o21a_1
XFILLER_0_136_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11901__B _03678_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08377_ _00429_ _00430_ _03982_ VGND VGND VPWR VPWR _00433_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_135_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12285__A _04714_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08482__B _00547_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07328_ net32 VGND VGND VPWR VPWR _02960_ sky130_fd_sc_hd__buf_4
XANTENNA__07379__A _03510_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07259_ _02072_ net184 VGND VGND VPWR VPWR _02204_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09594__A _03510_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10270_ _02311_ _02320_ _02503_ VGND VGND VPWR VPWR _02504_ sky130_fd_sc_hd__a21o_1
XANTENNA__07826__B net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11381__A1 _01312_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09326__A1 _00526_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13960_ _06541_ _06542_ VGND VGND VPWR VPWR _06543_ sky130_fd_sc_hd__nand2_1
X_12911_ _05363_ _05405_ VGND VGND VPWR VPWR _05407_ sky130_fd_sc_hd__and2_1
X_13891_ _06456_ _06466_ VGND VGND VPWR VPWR _06467_ sky130_fd_sc_hd__nor2_1
XANTENNA__11364__A _01312_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12842_ _05329_ _05330_ VGND VGND VPWR VPWR _05331_ sky130_fd_sc_hd__xnor2_1
XTAP_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12633__A1 _00392_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_632 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12773_ _05251_ _05253_ VGND VGND VPWR VPWR _05255_ sky130_fd_sc_hd__or2_1
XTAP_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12633__B2 _00389_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11724_ _04091_ _04100_ VGND VGND VPWR VPWR _04101_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09769__A _01955_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08673__A _02029_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_490 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11655_ _03889_ _04003_ VGND VGND VPWR VPWR _04025_ sky130_fd_sc_hd__xnor2_4
XANTENNA__11811__B _03748_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09488__B _00898_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07289__A net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10606_ _02870_ _02871_ VGND VGND VPWR VPWR _02873_ sky130_fd_sc_hd__xnor2_1
X_11586_ _03880_ _03948_ VGND VGND VPWR VPWR _03950_ sky130_fd_sc_hd__and2_1
XANTENNA__09262__B1 _01400_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07812__A1 _00563_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10537_ _03004_ _00293_ _02724_ _02728_ VGND VGND VPWR VPWR _02797_ sky130_fd_sc_hd__and4_1
X_13325_ _05844_ _05744_ _05845_ VGND VGND VPWR VPWR _05846_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_122_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07812__B2 _00639_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13256_ _05768_ _05779_ VGND VGND VPWR VPWR _05781_ sky130_fd_sc_hd__and2_1
X_10468_ _02720_ VGND VGND VPWR VPWR _02721_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__09935__C net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12207_ _04630_ _03682_ _00379_ _04632_ VGND VGND VPWR VPWR _04633_ sky130_fd_sc_hd__and4b_1
XANTENNA__07736__B net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13187_ _05705_ _05706_ _05710_ VGND VGND VPWR VPWR _05711_ sky130_fd_sc_hd__o21ai_4
X_10399_ _02121_ VGND VGND VPWR VPWR _02646_ sky130_fd_sc_hd__inv_2
XANTENNA__10175__A2 _03685_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12138_ _04481_ _04556_ VGND VGND VPWR VPWR _04557_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09009__A _03004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12069_ _03929_ _04480_ VGND VGND VPWR VPWR _04481_ sky130_fd_sc_hd__nor2_1
XANTENNA__08848__A _05577_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09868__A2 _00755_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09219__B_N _01352_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08540__A2 _04026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08300_ _04334_ _00348_ VGND VGND VPWR VPWR _00349_ sky130_fd_sc_hd__xor2_2
XFILLER_0_87_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09280_ _01409_ _01420_ VGND VGND VPWR VPWR _01421_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08231_ _05566_ _06775_ VGND VGND VPWR VPWR _00275_ sky130_fd_sc_hd__nand2_1
XFILLER_0_118_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09398__B net49 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08162_ _00204_ _00205_ VGND VGND VPWR VPWR _00206_ sky130_fd_sc_hd__or2_4
XFILLER_0_132_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07113_ _00584_ _00595_ VGND VGND VPWR VPWR _00606_ sky130_fd_sc_hd__and2b_1
X_08093_ _00134_ _00136_ VGND VGND VPWR VPWR _00137_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11449__A _00262_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08995_ _01062_ VGND VGND VPWR VPWR _01108_ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09587__A2_N _01486_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07946_ _07041_ _07074_ VGND VGND VPWR VPWR _07075_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_98_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07877_ _06951_ _06971_ VGND VGND VPWR VPWR _07006_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08531__A2 _00376_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09616_ _01605_ _01786_ VGND VGND VPWR VPWR _01789_ sky130_fd_sc_hd__or2_1
XFILLER_0_92_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09547_ _01697_ _01712_ VGND VGND VPWR VPWR _01713_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_78_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09478_ _01056_ _01238_ _01243_ VGND VGND VPWR VPWR _01638_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_136_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08429_ _00487_ _00489_ VGND VGND VPWR VPWR _00490_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09739__D net52 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11440_ _03757_ _03782_ _03788_ VGND VGND VPWR VPWR _03789_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_135_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire137 _06364_ VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__buf_1
XFILLER_0_104_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11371_ _03690_ _03689_ _03688_ VGND VGND VPWR VPWR _03713_ sky130_fd_sc_hd__a21bo_1
XANTENNA__13591__A2 _02856_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10322_ _02214_ _02546_ _02547_ _02560_ VGND VGND VPWR VPWR _02561_ sky130_fd_sc_hd__and4_1
X_13110_ _05154_ _05625_ _05218_ VGND VGND VPWR VPWR _05626_ sky130_fd_sc_hd__o21a_2
XANTENNA__07837__A _06875_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14090_ _05960_ _06619_ VGND VGND VPWR VPWR _06685_ sky130_fd_sc_hd__nor2_1
XFILLER_0_131_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13041_ _04604_ VGND VGND VPWR VPWR _05550_ sky130_fd_sc_hd__inv_2
X_10253_ _02242_ _02269_ _02151_ VGND VGND VPWR VPWR _02486_ sky130_fd_sc_hd__a21oi_2
XANTENNA__11354__A1 _02246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11354__B2 _02249_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12551__B1 _01289_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10184_ _02399_ _02409_ VGND VGND VPWR VPWR _02410_ sky130_fd_sc_hd__xor2_2
XFILLER_0_100_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12303__B1 _02189_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13943_ _06331_ _06355_ VGND VGND VPWR VPWR _06524_ sky130_fd_sc_hd__xor2_2
XFILLER_0_88_316 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13874_ _06442_ _06444_ VGND VGND VPWR VPWR _06448_ sky130_fd_sc_hd__nor2_1
XFILLER_0_69_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12825_ _05140_ _05218_ _05311_ VGND VGND VPWR VPWR _05312_ sky130_fd_sc_hd__a21o_1
XFILLER_0_29_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12918__A _01108_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12756_ _00607_ _03738_ VGND VGND VPWR VPWR _05237_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11707_ _04061_ _04082_ VGND VGND VPWR VPWR _04083_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12687_ _05080_ _05160_ VGND VGND VPWR VPWR _05161_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09011__B _00151_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11638_ _03868_ _03874_ _03871_ VGND VGND VPWR VPWR _04007_ sky130_fd_sc_hd__and3_1
XFILLER_0_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11569_ _03919_ _03921_ VGND VGND VPWR VPWR _03931_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_25_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07169__D _01208_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07747__A _01383_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13308_ _05819_ _05826_ _05829_ VGND VGND VPWR VPWR _05830_ sky130_fd_sc_hd__a21o_1
XFILLER_0_122_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09665__C _00145_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12372__B _00457_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13239_ _01640_ _02046_ _02492_ _05763_ VGND VGND VPWR VPWR _05765_ sky130_fd_sc_hd__nand4_2
XFILLER_0_0_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07800_ _06911_ _06928_ VGND VGND VPWR VPWR _06929_ sky130_fd_sc_hd__xor2_2
X_08780_ _00841_ _00873_ VGND VGND VPWR VPWR _00874_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_46_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07731_ _02664_ _00475_ VGND VGND VPWR VPWR _06860_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08513__A2 _03894_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07662_ _06604_ _06340_ VGND VGND VPWR VPWR _06615_ sky130_fd_sc_hd__xnor2_1
X_09401_ _01419_ _01551_ VGND VGND VPWR VPWR _01553_ sky130_fd_sc_hd__nor2_1
X_07593_ _05837_ _05847_ VGND VGND VPWR VPWR _05857_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09332_ _01315_ _01475_ VGND VGND VPWR VPWR _01477_ sky130_fd_sc_hd__and2_1
XFILLER_0_87_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09263_ _01066_ _01399_ _01401_ VGND VGND VPWR VPWR _01402_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_63_706 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11451__B _00121_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09559__D _01472_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08214_ _00114_ VGND VGND VPWR VPWR _00258_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_118_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09226__B1 _00380_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09194_ _01324_ _01325_ VGND VGND VPWR VPWR _01326_ sky130_fd_sc_hd__and2b_1
XFILLER_0_117_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08145_ _00186_ _00188_ _00183_ VGND VGND VPWR VPWR _00189_ sky130_fd_sc_hd__and3_1
XFILLER_0_126_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08076_ _00021_ _00022_ _00023_ VGND VGND VPWR VPWR _00120_ sky130_fd_sc_hd__and3_1
XANTENNA__13378__B _01505_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13809__D _03686_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09591__B _06820_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13711__A2_N _02721_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08978_ _01088_ _01089_ VGND VGND VPWR VPWR _01090_ sky130_fd_sc_hd__and2b_1
X_07929_ _00672_ _05027_ _06901_ _06900_ VGND VGND VPWR VPWR _07058_ sky130_fd_sc_hd__a31o_1
XANTENNA__07823__C net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10940_ _03199_ _03204_ _03192_ VGND VGND VPWR VPWR _03240_ sky130_fd_sc_hd__o21a_1
XANTENNA__10311__A2 _01368_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08000__B _02040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10871_ _03159_ _03161_ _03163_ VGND VGND VPWR VPWR _03164_ sky130_fd_sc_hd__o21a_1
X_12610_ _05074_ _05075_ VGND VGND VPWR VPWR _05076_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_66_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13261__A1 _02278_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13590_ _01181_ _01250_ _02856_ _02858_ VGND VGND VPWR VPWR _06136_ sky130_fd_sc_hd__and4_1
XFILLER_0_38_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11361__B _00844_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12541_ _04864_ _04865_ VGND VGND VPWR VPWR _05000_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_54_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13013__A1 _05509_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12472_ _04919_ _04920_ VGND VGND VPWR VPWR _04924_ sky130_fd_sc_hd__nor2_1
XANTENNA__08951__A _01059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14211_ _06800_ VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11423_ _03736_ _03739_ _03746_ VGND VGND VPWR VPWR _03770_ sky130_fd_sc_hd__or3_1
XFILLER_0_105_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14142_ _06736_ _06739_ VGND VGND VPWR VPWR _06740_ sky130_fd_sc_hd__and2b_1
X_11354_ _02246_ _01957_ _03690_ _02249_ VGND VGND VPWR VPWR _03694_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_21_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07567__A _05577_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10305_ _02502_ _02541_ VGND VGND VPWR VPWR _02542_ sky130_fd_sc_hd__xnor2_1
X_14073_ _06664_ _06665_ VGND VGND VPWR VPWR _06666_ sky130_fd_sc_hd__or2_1
X_11285_ _03617_ _03608_ _03618_ VGND VGND VPWR VPWR _03619_ sky130_fd_sc_hd__o21ai_1
XTAP_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13024_ _05512_ _05514_ _05515_ _05513_ VGND VGND VPWR VPWR _05531_ sky130_fd_sc_hd__a22o_1
X_10236_ _02139_ _02465_ VGND VGND VPWR VPWR _02468_ sky130_fd_sc_hd__nand2_1
X_10167_ _02074_ _02080_ _02075_ VGND VGND VPWR VPWR _02392_ sky130_fd_sc_hd__a21bo_1
XANTENNA__11536__B _06874_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10098_ _04081_ net53 VGND VGND VPWR VPWR _02316_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13926_ _06491_ _06493_ _06501_ _06503_ VGND VGND VPWR VPWR _06506_ sky130_fd_sc_hd__o22a_1
XFILLER_0_89_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13857_ _05918_ _06426_ _06429_ VGND VGND VPWR VPWR _06430_ sky130_fd_sc_hd__and3_1
XFILLER_0_76_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08845__B _00639_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12808_ _05292_ _05293_ VGND VGND VPWR VPWR _05294_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13788_ _06341_ _06342_ _06335_ _06338_ VGND VGND VPWR VPWR _06354_ sky130_fd_sc_hd__o211a_1
XFILLER_0_29_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12739_ _05155_ _05216_ _05217_ VGND VGND VPWR VPWR _05218_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_32_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08283__D _06874_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08861__A _01372_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_142_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_822 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09950_ _01921_ _01926_ VGND VGND VPWR VPWR _02154_ sky130_fd_sc_hd__nand2_1
XANTENNA__07196__B _00978_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07627__D _03268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08901_ _00813_ _01004_ VGND VGND VPWR VPWR _01006_ sky130_fd_sc_hd__and2_1
XFILLER_0_110_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09881_ _03521_ _00486_ _00413_ _00572_ VGND VGND VPWR VPWR _02078_ sky130_fd_sc_hd__and4_1
XANTENNA__11869__A2 _01600_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08832_ _00758_ _00928_ VGND VGND VPWR VPWR _00930_ sky130_fd_sc_hd__and2b_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14103__A _06684_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08763_ _00484_ _00490_ _00684_ VGND VGND VPWR VPWR _00855_ sky130_fd_sc_hd__o21a_1
XANTENNA__08101__A _00144_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07714_ _06831_ _06830_ VGND VGND VPWR VPWR _06843_ sky130_fd_sc_hd__and2b_1
XFILLER_0_79_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12294__A2 _02426_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08694_ _00778_ VGND VGND VPWR VPWR _00779_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_68_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07645_ _06417_ VGND VGND VPWR VPWR _06428_ sky130_fd_sc_hd__buf_4
XFILLER_0_95_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08755__B _00843_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07576_ _05511_ net190 VGND VGND VPWR VPWR _05687_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_48_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11181__B _03480_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09315_ _00262_ _00859_ _01136_ VGND VGND VPWR VPWR _01458_ sky130_fd_sc_hd__and3_1
XFILLER_0_118_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09246_ _03268_ _00612_ _00613_ _05577_ VGND VGND VPWR VPWR _01384_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_35_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08670__A1 _05731_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08670__B2 _01000_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_435 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09586__B _01486_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09177_ _01245_ _01305_ VGND VGND VPWR VPWR _01308_ sky130_fd_sc_hd__and2_1
XFILLER_0_90_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12293__A _00575_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_411 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_496 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08128_ _00170_ _00171_ VGND VGND VPWR VPWR _00172_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_71_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12754__B1 _01254_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08059_ _00102_ VGND VGND VPWR VPWR _00103_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10780__A2 _02720_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11070_ _03373_ _03381_ _03382_ VGND VGND VPWR VPWR _03383_ sky130_fd_sc_hd__a21oi_1
Xoutput68 net68 VGND VGND VPWR VPWR prod[12] sky130_fd_sc_hd__clkbuf_4
Xoutput79 net79 VGND VGND VPWR VPWR prod[22] sky130_fd_sc_hd__clkbuf_4
X_10021_ _02228_ _02231_ VGND VGND VPWR VPWR _02232_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11972_ _04308_ _04310_ _04373_ VGND VGND VPWR VPWR _04374_ sky130_fd_sc_hd__and3_1
XANTENNA__08946__A _00898_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13711_ _02427_ _02721_ _06254_ _06255_ VGND VGND VPWR VPWR _06269_ sky130_fd_sc_hd__o2bb2a_1
X_10923_ _03207_ _03220_ VGND VGND VPWR VPWR _03221_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_86_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11372__A _01155_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13642_ _05978_ _06192_ VGND VGND VPWR VPWR _06193_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10854_ _03141_ _03144_ VGND VGND VPWR VPWR _03145_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13573_ _05978_ _05991_ VGND VGND VPWR VPWR _06117_ sky130_fd_sc_hd__and2_1
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10785_ _03064_ _03067_ VGND VGND VPWR VPWR _03069_ sky130_fd_sc_hd__or2_1
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_834 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11796__A1 _01361_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11796__B2 _01405_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12524_ _04941_ _04943_ _04938_ VGND VGND VPWR VPWR _04981_ sky130_fd_sc_hd__a21bo_1
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09777__A _01295_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12455_ _04903_ _04904_ VGND VGND VPWR VPWR _04905_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11548__A1 _06964_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11548__B2 _00121_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11406_ _00257_ _00670_ _03750_ _03748_ VGND VGND VPWR VPWR _03752_ sky130_fd_sc_hd__nand4_1
XFILLER_0_1_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07728__C net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12386_ _00782_ _00613_ _00571_ _00734_ VGND VGND VPWR VPWR _04830_ sky130_fd_sc_hd__and4_1
X_14125_ _06720_ _06721_ VGND VGND VPWR VPWR _06722_ sky130_fd_sc_hd__nor2_1
XANTENNA__08964__A2 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11337_ _03638_ _03665_ _03627_ VGND VGND VPWR VPWR _03676_ sky130_fd_sc_hd__a21o_1
XANTENNA_output77_A net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14056_ _06610_ _06647_ VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__xnor2_4
X_11268_ _03599_ _03600_ VGND VGND VPWR VPWR _03601_ sky130_fd_sc_hd__and2_1
XFILLER_0_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13007_ _04575_ _04580_ _04584_ VGND VGND VPWR VPWR _05513_ sky130_fd_sc_hd__o21ai_4
XANTENNA__11547__A _06965_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10219_ _02448_ VGND VGND VPWR VPWR _02449_ sky130_fd_sc_hd__inv_2
X_11199_ _03388_ _03396_ _03401_ VGND VGND VPWR VPWR _03525_ sky130_fd_sc_hd__nor3_1
XFILLER_0_89_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13481__B _01415_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13909_ _06365_ _06376_ _06414_ _06486_ VGND VGND VPWR VPWR _06487_ sky130_fd_sc_hd__nor4_1
XFILLER_0_49_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07430_ _01284_ VGND VGND VPWR VPWR _04081_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_147_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07361_ _03279_ _03312_ VGND VGND VPWR VPWR _03323_ sky130_fd_sc_hd__xor2_1
XFILLER_0_45_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09100_ _00932_ _01190_ _01223_ VGND VGND VPWR VPWR _01224_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_45_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07292_ net60 net26 VGND VGND VPWR VPWR _02565_ sky130_fd_sc_hd__nand2_1
XANTENNA__07455__A2 _00388_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_142_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09031_ _01147_ VGND VGND VPWR VPWR _01148_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12841__A _00745_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09933_ _02134_ VGND VGND VPWR VPWR _02135_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09864_ _00004_ _00390_ _00393_ _07004_ VGND VGND VPWR VPWR _02059_ sky130_fd_sc_hd__a22o_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09380__A2 _00605_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08815_ _00738_ _00909_ VGND VGND VPWR VPWR _00911_ sky130_fd_sc_hd__and2_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09795_ _05456_ _00138_ _00572_ _01586_ VGND VGND VPWR VPWR _01984_ sky130_fd_sc_hd__and4_1
XFILLER_0_84_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08746_ _00816_ _00835_ VGND VGND VPWR VPWR _00837_ sky130_fd_sc_hd__xor2_1
XTAP_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08766__A _00310_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10278__A1 _01372_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13391__B _01517_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08677_ _00758_ _00760_ VGND VGND VPWR VPWR _00761_ sky130_fd_sc_hd__or2_2
XFILLER_0_95_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07628_ _02007_ _05566_ _06197_ _06219_ VGND VGND VPWR VPWR _06241_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_95_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07694__A2 _06818_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07559_ _05456_ _01350_ _05489_ VGND VGND VPWR VPWR _05500_ sky130_fd_sc_hd__and3_1
XFILLER_0_48_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_536 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_845 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10570_ _02816_ _02832_ VGND VGND VPWR VPWR _02833_ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09597__A _00475_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07446__A2 net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09229_ _01362_ _01364_ VGND VGND VPWR VPWR _01365_ sky130_fd_sc_hd__or2_1
XFILLER_0_118_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07829__B _06744_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_243 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12240_ _04654_ _04655_ _04652_ VGND VGND VPWR VPWR _04669_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_133_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12171_ _04545_ _04592_ _04539_ VGND VGND VPWR VPWR _04593_ sky130_fd_sc_hd__o21ai_1
XANTENNA__13847__A _02189_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10753__A2 _02765_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11122_ _03412_ _03417_ _03404_ VGND VGND VPWR VPWR _03440_ sky130_fd_sc_hd__o21a_1
XFILLER_0_102_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11053_ _03342_ _03344_ _03363_ _03339_ VGND VGND VPWR VPWR _03364_ sky130_fd_sc_hd__a211o_1
X_10004_ _04598_ _00612_ _00613_ _05192_ VGND VGND VPWR VPWR _02213_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11955_ _04122_ _04141_ _04285_ _04254_ VGND VGND VPWR VPWR _04355_ sky130_fd_sc_hd__a211o_1
XANTENNA_output115_A net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10906_ _03197_ _03198_ VGND VGND VPWR VPWR _03203_ sky130_fd_sc_hd__and2_1
XFILLER_0_80_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11886_ _04272_ _04277_ VGND VGND VPWR VPWR _04280_ sky130_fd_sc_hd__nand2_1
X_13625_ _06008_ _06047_ VGND VGND VPWR VPWR _06174_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10837_ _02512_ _02515_ _03126_ VGND VGND VPWR VPWR _03127_ sky130_fd_sc_hd__a21o_1
XFILLER_0_67_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11769__A1 _02007_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11769__B2 _01178_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13556_ _06091_ _06097_ VGND VGND VPWR VPWR _06099_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10768_ _03003_ _03050_ VGND VGND VPWR VPWR _03051_ sky130_fd_sc_hd__nor2_1
XFILLER_0_125_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12507_ _04059_ _03938_ VGND VGND VPWR VPWR _04963_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07739__B _06744_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13487_ _01415_ _03697_ VGND VGND VPWR VPWR _06023_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10699_ _02973_ _02974_ VGND VGND VPWR VPWR _02975_ sky130_fd_sc_hd__nand2_1
XFILLER_0_124_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12438_ _04827_ _04875_ VGND VGND VPWR VPWR _04887_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_2_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12369_ _04809_ _04810_ VGND VGND VPWR VPWR _04811_ sky130_fd_sc_hd__nand2_1
X_14108_ _06078_ _02743_ _04014_ _02742_ VGND VGND VPWR VPWR _06704_ sky130_fd_sc_hd__and4_1
XANTENNA__07755__A _02259_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14039_ net135 _06629_ _06578_ VGND VGND VPWR VPWR _06630_ sky130_fd_sc_hd__or3_2
XFILLER_0_38_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11427__D _01249_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08600_ _00479_ _00675_ VGND VGND VPWR VPWR _00677_ sky130_fd_sc_hd__nor2_1
XANTENNA__08570__B1 _00151_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09580_ _01465_ _01723_ _01748_ VGND VGND VPWR VPWR _01749_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_54_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07490__A net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08531_ _02259_ _00376_ _00379_ _02171_ VGND VGND VPWR VPWR _00601_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_77_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07125__A1 net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07125__B2 _00573_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08462_ _07040_ VGND VGND VPWR VPWR _00526_ sky130_fd_sc_hd__buf_4
XANTENNA__11443__C _02133_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07413_ net10 VGND VGND VPWR VPWR _03894_ sky130_fd_sc_hd__clkbuf_4
X_08393_ _00444_ _00449_ VGND VGND VPWR VPWR _00450_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_856 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07344_ net60 net26 _02543_ _02532_ VGND VGND VPWR VPWR _03136_ sky130_fd_sc_hd__a31o_1
XFILLER_0_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07275_ _02193_ _02368_ VGND VGND VPWR VPWR _02379_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_60_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09014_ _01119_ _01121_ _01128_ VGND VGND VPWR VPWR _01129_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_5_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_596 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13667__A _01108_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07665__A _06626_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09916_ _01564_ VGND VGND VPWR VPWR _02117_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__10091__A _01350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09847_ _01828_ _01759_ VGND VGND VPWR VPWR _02042_ sky130_fd_sc_hd__or2_1
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11696__B1 _01211_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09778_ _01306_ net19 VGND VGND VPWR VPWR _01966_ sky130_fd_sc_hd__nand2_1
XTAP_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08729_ _00294_ VGND VGND VPWR VPWR _00818_ sky130_fd_sc_hd__clkbuf_4
XTAP_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ _04039_ _04118_ VGND VGND VPWR VPWR _04119_ sky130_fd_sc_hd__nor2_1
XANTENNA__11353__C _01956_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10671__A1 _05181_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10671__B2 _00094_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11671_ _07010_ _00423_ _03762_ _00101_ VGND VGND VPWR VPWR _04043_ sky130_fd_sc_hd__a22oi_1
XTAP_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13410_ _05248_ _05399_ _05400_ _01956_ _04714_ VGND VGND VPWR VPWR _05939_ sky130_fd_sc_hd__a32o_1
XFILLER_0_64_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10622_ _02887_ _02889_ VGND VGND VPWR VPWR _02890_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_675 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10423__A1 _00311_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13341_ _05862_ _05860_ VGND VGND VPWR VPWR _05863_ sky130_fd_sc_hd__nor2_1
XANTENNA__07559__B _01350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10553_ _00377_ _02993_ _02168_ _02723_ VGND VGND VPWR VPWR _02814_ sky130_fd_sc_hd__and4_1
XFILLER_0_106_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13272_ _05474_ _05490_ VGND VGND VPWR VPWR _05796_ sky130_fd_sc_hd__and2_1
X_10484_ _01473_ _02247_ _02736_ _02737_ VGND VGND VPWR VPWR _02738_ sky130_fd_sc_hd__nand4_1
XFILLER_0_20_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12223_ _00778_ _01248_ _02117_ _00783_ VGND VGND VPWR VPWR _04650_ sky130_fd_sc_hd__a22o_1
XANTENNA__13577__A _01249_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09774__B _01960_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12154_ _04562_ _04564_ _04557_ VGND VGND VPWR VPWR _04574_ sky130_fd_sc_hd__o21a_1
XANTENNA__09592__A2 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11105_ _03416_ _03420_ VGND VGND VPWR VPWR _03421_ sky130_fd_sc_hd__xnor2_1
X_12085_ _04496_ _04416_ _04419_ VGND VGND VPWR VPWR _04498_ sky130_fd_sc_hd__nor3_1
X_11036_ _00142_ _04037_ _02566_ _02564_ _00778_ VGND VGND VPWR VPWR _03346_ sky130_fd_sc_hd__a32o_1
XANTENNA__14201__A _00344_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12987_ _05474_ _05490_ VGND VGND VPWR VPWR _05491_ sky130_fd_sc_hd__xor2_1
XFILLER_0_86_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11938_ _04258_ _04260_ _04336_ VGND VGND VPWR VPWR _04337_ sky130_fd_sc_hd__o21a_1
XFILLER_0_115_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11869_ _06775_ _01600_ _04034_ _04033_ _00575_ VGND VGND VPWR VPWR _04261_ sky130_fd_sc_hd__a32o_1
XFILLER_0_55_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13608_ _06154_ _06155_ VGND VGND VPWR VPWR _06156_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_145_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13539_ _06075_ _06077_ _06078_ _06074_ VGND VGND VPWR VPWR _06080_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_40_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14156__A2 _05833_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13487__A _01415_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13364__B1 _02721_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12391__A _01518_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07485__A net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11719__B _01585_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07962_ _02259_ _02171_ _00004_ _06885_ VGND VGND VPWR VPWR _00006_ sky130_fd_sc_hd__and4_1
X_09701_ _01870_ _01871_ _01879_ VGND VGND VPWR VPWR _01881_ sky130_fd_sc_hd__or3_1
XFILLER_0_4_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07346__A1 _01044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07893_ _00639_ _06818_ _06820_ net29 VGND VGND VPWR VPWR _07022_ sky130_fd_sc_hd__a22oi_1
XANTENNA__08543__B1 _00613_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09632_ _01803_ _01805_ VGND VGND VPWR VPWR _01806_ sky130_fd_sc_hd__xnor2_2
XANTENNA__13419__A1 _01183_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13419__B2 _01108_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09563_ _00544_ _00859_ _01728_ VGND VGND VPWR VPWR _01730_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_77_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08514_ _01361_ _01405_ _03773_ _03938_ VGND VGND VPWR VPWR _00582_ sky130_fd_sc_hd__nand4_1
XFILLER_0_38_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09494_ _01652_ _01653_ VGND VGND VPWR VPWR _01654_ sky130_fd_sc_hd__xor2_1
XANTENNA__08846__A1 _05742_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08846__B2 _00563_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08445_ _00505_ _00506_ VGND VGND VPWR VPWR _00507_ sky130_fd_sc_hd__nor2_1
XFILLER_0_65_428 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08376_ _03982_ _00429_ _00430_ VGND VGND VPWR VPWR _00432_ sky130_fd_sc_hd__and3_1
XFILLER_0_147_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12285__B _01181_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07327_ _00344_ _00410_ _02927_ _02938_ VGND VGND VPWR VPWR _02949_ sky130_fd_sc_hd__a31o_1
XFILLER_0_144_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07258_ _00683_ _02182_ VGND VGND VPWR VPWR _02193_ sky130_fd_sc_hd__or2_1
XFILLER_0_60_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07189_ _01328_ _01427_ VGND VGND VPWR VPWR _01438_ sky130_fd_sc_hd__and2_1
XANTENNA__09023__A1 _03543_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09594__B _03762_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07395__A _03685_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12910_ _05363_ _05405_ VGND VGND VPWR VPWR _05406_ sky130_fd_sc_hd__nor2_1
X_13890_ _06454_ _06455_ VGND VGND VPWR VPWR _06466_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11364__B _03680_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12841_ _00745_ _02168_ VGND VGND VPWR VPWR _05330_ sky130_fd_sc_hd__nand2_1
XTAP_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12772_ _05251_ _05253_ VGND VGND VPWR VPWR _05254_ sky130_fd_sc_hd__and2_1
XTAP_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12633__A2 _02168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_644 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ _04098_ _04099_ VGND VGND VPWR VPWR _04100_ sky130_fd_sc_hd__nor2_1
XTAP_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08673__B _00755_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11654_ _04023_ VGND VGND VPWR VPWR _04024_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_804 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10605_ _00144_ _01412_ VGND VGND VPWR VPWR _02871_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09262__A1 _02171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07289__B net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11585_ _03878_ _03879_ VGND VGND VPWR VPWR _03948_ sky130_fd_sc_hd__or2_1
XANTENNA__09262__B2 _02467_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13324_ _05748_ _05646_ VGND VGND VPWR VPWR _05845_ sky130_fd_sc_hd__nor2_1
X_10536_ _02770_ _02794_ VGND VGND VPWR VPWR _02796_ sky130_fd_sc_hd__nand2_2
XANTENNA__07812__A2 _06818_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13255_ _05524_ _05546_ VGND VGND VPWR VPWR _05779_ sky130_fd_sc_hd__and2_1
X_10467_ _02169_ VGND VGND VPWR VPWR _02720_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_110_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09935__D _02133_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12206_ _00784_ _01953_ _02134_ _00374_ VGND VGND VPWR VPWR _04632_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13186_ _05705_ _05706_ _05708_ VGND VGND VPWR VPWR _05710_ sky130_fd_sc_hd__a21o_1
X_10398_ _02596_ _02644_ VGND VGND VPWR VPWR _02645_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__07736__C net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12137_ _04482_ _04479_ VGND VGND VPWR VPWR _04556_ sky130_fd_sc_hd__and2b_1
XANTENNA__09009__B _00113_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10580__B1 _02305_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12068_ _03554_ _01183_ _01252_ _00530_ VGND VGND VPWR VPWR _04480_ sky130_fd_sc_hd__a22oi_1
XANTENNA__08848__B _04026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11019_ _03324_ _03325_ VGND VGND VPWR VPWR _03327_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08864__A _01230_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12386__A _00782_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08230_ _00102_ _00105_ VGND VGND VPWR VPWR _00274_ sky130_fd_sc_hd__or2_1
XFILLER_0_74_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10618__B _04939_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08161_ _06998_ _00203_ _00202_ VGND VGND VPWR VPWR _00205_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_16_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09695__A _02960_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07112_ _00563_ _00573_ net44 net28 VGND VGND VPWR VPWR _00595_ sky130_fd_sc_hd__a22o_1
XFILLER_0_113_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08092_ _07003_ _07036_ _00040_ _00135_ VGND VGND VPWR VPWR _00136_ sky130_fd_sc_hd__a31o_1
XFILLER_0_70_442 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14106__A _02743_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11449__B _03680_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12560__A1 _00390_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08994_ _00464_ _01062_ _01106_ VGND VGND VPWR VPWR _01107_ sky130_fd_sc_hd__and3_1
X_07945_ _07073_ _07072_ VGND VGND VPWR VPWR _07074_ sky130_fd_sc_hd__and2b_1
X_07876_ _02467_ _07004_ VGND VGND VPWR VPWR _07005_ sky130_fd_sc_hd__nand2_1
X_09615_ _01605_ _01786_ VGND VGND VPWR VPWR _01787_ sky130_fd_sc_hd__nand2_1
X_09546_ _01709_ _01710_ VGND VGND VPWR VPWR _01712_ sky130_fd_sc_hd__or2_2
XFILLER_0_66_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09477_ _01239_ VGND VGND VPWR VPWR _01637_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08428_ _00255_ _00266_ _00488_ VGND VGND VPWR VPWR _00489_ sky130_fd_sc_hd__a21o_1
XFILLER_0_18_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08359_ net13 VGND VGND VPWR VPWR _00413_ sky130_fd_sc_hd__buf_2
XFILLER_0_61_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_656 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11370_ _03692_ net142 _03710_ VGND VGND VPWR VPWR _03712_ sky130_fd_sc_hd__nor3_1
XFILLER_0_116_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10321_ _02558_ _02559_ VGND VGND VPWR VPWR _02560_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13040_ _05536_ _05538_ VGND VGND VPWR VPWR _05549_ sky130_fd_sc_hd__xor2_2
X_10252_ _02242_ _02269_ VGND VGND VPWR VPWR _02485_ sky130_fd_sc_hd__nor2_1
XANTENNA__11354__A2 _01957_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12551__A1 _00376_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12551__B2 _00380_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10183_ _02407_ _02408_ VGND VGND VPWR VPWR _02409_ sky130_fd_sc_hd__nand2_2
XANTENNA__08949__A net49 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12303__A1 _01288_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12303__B2 _00416_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13942_ _06508_ _06522_ VGND VGND VPWR VPWR _06523_ sky130_fd_sc_hd__nor2_1
X_13873_ _06401_ _06446_ VGND VGND VPWR VPWR _06447_ sky130_fd_sc_hd__and2_1
XFILLER_0_88_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13590__A _01181_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12824_ _05307_ _05310_ VGND VGND VPWR VPWR _05311_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12918__B _01183_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12755_ _01180_ _05233_ _05234_ VGND VGND VPWR VPWR _05235_ sky130_fd_sc_hd__a21bo_1
XTAP_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11706_ _04075_ _04080_ VGND VGND VPWR VPWR _04082_ sky130_fd_sc_hd__xor2_1
XFILLER_0_56_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12686_ _05078_ _05079_ VGND VGND VPWR VPWR _05160_ sky130_fd_sc_hd__and2_1
XFILLER_0_71_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11637_ _03889_ _04003_ _04005_ VGND VGND VPWR VPWR _04006_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_25_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07246__B1 _02040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11568_ _03928_ _03929_ VGND VGND VPWR VPWR _03930_ sky130_fd_sc_hd__and2b_1
XFILLER_0_80_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13307_ _05745_ _05738_ _05828_ VGND VGND VPWR VPWR _05829_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_122_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10519_ _02775_ _02776_ VGND VGND VPWR VPWR _02777_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10454__A _02482_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07747__B _06875_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11499_ _03717_ _03720_ VGND VGND VPWR VPWR _03854_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09665__D _04917_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13238_ _02494_ _05763_ VGND VGND VPWR VPWR _05764_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13169_ _05196_ _05206_ VGND VGND VPWR VPWR _05691_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_137_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07730_ _06857_ _06858_ VGND VGND VPWR VPWR _06859_ sky130_fd_sc_hd__and2b_1
XFILLER_0_46_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09171__B1 _00393_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07661_ _06582_ _06593_ VGND VGND VPWR VPWR _06604_ sky130_fd_sc_hd__nor2_1
X_09400_ _01419_ _01551_ VGND VGND VPWR VPWR _01552_ sky130_fd_sc_hd__and2_1
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07592_ _02007_ _05588_ VGND VGND VPWR VPWR _05847_ sky130_fd_sc_hd__nand2_1
XANTENNA__08594__A _00258_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09331_ _01315_ _01475_ VGND VGND VPWR VPWR _01476_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10629__A _00819_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09262_ _02171_ _00460_ _01400_ _02467_ VGND VGND VPWR VPWR _01401_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11451__C _01953_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08213_ _00113_ VGND VGND VPWR VPWR _00257_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_90_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09226__A1 _00410_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09193_ _01018_ _01132_ _01129_ VGND VGND VPWR VPWR _01325_ sky130_fd_sc_hd__o21a_1
XFILLER_0_133_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09226__B2 _03015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_431 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08144_ _07000_ _00187_ VGND VGND VPWR VPWR _00188_ sky130_fd_sc_hd__nor2_1
XANTENNA__07788__A1 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12781__A1 _02305_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08075_ _00117_ _00118_ VGND VGND VPWR VPWR _00119_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_113_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_648 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07673__A net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08977_ _00541_ _04103_ _04191_ _00639_ VGND VGND VPWR VPWR _01089_ sky130_fd_sc_hd__a22o_1
XANTENNA__09591__C net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07928_ _06904_ _06907_ _07056_ VGND VGND VPWR VPWR _07057_ sky130_fd_sc_hd__a21bo_1
XANTENNA__07823__D net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07859_ _05368_ _05390_ VGND VGND VPWR VPWR _06988_ sky130_fd_sc_hd__and2_1
XANTENNA__08000__C _04917_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10870_ _03154_ _03162_ VGND VGND VPWR VPWR _03163_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09529_ _01540_ VGND VGND VPWR VPWR _01693_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12540_ _04944_ _04979_ VGND VGND VPWR VPWR _04999_ sky130_fd_sc_hd__xor2_2
XFILLER_0_109_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11361__C _03687_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12471_ _04766_ _04922_ VGND VGND VPWR VPWR _04923_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14210_ _01766_ _06799_ VGND VGND VPWR VPWR _06800_ sky130_fd_sc_hd__and2_1
XFILLER_0_124_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11422_ _07004_ _03748_ _03763_ _03768_ VGND VGND VPWR VPWR _03769_ sky130_fd_sc_hd__a31o_1
XFILLER_0_61_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14141_ _06673_ _06737_ _06738_ VGND VGND VPWR VPWR _06739_ sky130_fd_sc_hd__o21a_1
XFILLER_0_104_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11353_ _02246_ _02249_ _01956_ _03687_ VGND VGND VPWR VPWR _03693_ sky130_fd_sc_hd__and4_1
XFILLER_0_22_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10304_ _02538_ _02540_ VGND VGND VPWR VPWR _02541_ sky130_fd_sc_hd__xor2_2
X_14072_ _06662_ _06663_ _06077_ _04014_ VGND VGND VPWR VPWR _06665_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11284_ _03597_ _03601_ VGND VGND VPWR VPWR _03618_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13023_ _05509_ _05529_ VGND VGND VPWR VPWR _05530_ sky130_fd_sc_hd__xnor2_1
X_10235_ _02139_ _02465_ VGND VGND VPWR VPWR _02466_ sky130_fd_sc_hd__or2_1
X_10166_ _02145_ _02147_ VGND VGND VPWR VPWR _02391_ sky130_fd_sc_hd__or2b_1
X_10097_ _02312_ _02172_ _02314_ VGND VGND VPWR VPWR _02315_ sky130_fd_sc_hd__a21bo_1
XANTENNA__11536__C _01177_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13925_ _06491_ _06493_ _06501_ _06503_ VGND VGND VPWR VPWR _06504_ sky130_fd_sc_hd__nor4_1
XANTENNA__07703__A1 net149 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13856_ _05921_ _05926_ _06427_ VGND VGND VPWR VPWR _06429_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_76_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12807_ _05054_ _05289_ _05290_ _05288_ VGND VGND VPWR VPWR _05293_ sky130_fd_sc_hd__a31o_1
XFILLER_0_9_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13787_ _06348_ _06352_ VGND VGND VPWR VPWR _06353_ sky130_fd_sc_hd__nand2_1
X_10999_ _03303_ _03304_ VGND VGND VPWR VPWR _03305_ sky130_fd_sc_hd__nor2_2
XFILLER_0_146_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12738_ _05132_ _05139_ VGND VGND VPWR VPWR _05217_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12669_ _04896_ _04910_ _05035_ VGND VGND VPWR VPWR _05141_ sky130_fd_sc_hd__and3_1
XANTENNA__08861__B net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08900_ _00813_ _01004_ VGND VGND VPWR VPWR _01005_ sky130_fd_sc_hd__nor2_1
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09880_ _03554_ _00416_ _01288_ _00508_ VGND VGND VPWR VPWR _02077_ sky130_fd_sc_hd__a22o_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08831_ _00591_ _00757_ _00928_ VGND VGND VPWR VPWR _00929_ sky130_fd_sc_hd__nor3_1
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08762_ _00685_ VGND VGND VPWR VPWR _00854_ sky130_fd_sc_hd__inv_2
X_07713_ _00880_ net63 VGND VGND VPWR VPWR _06842_ sky130_fd_sc_hd__nand2_1
X_08693_ _00777_ VGND VGND VPWR VPWR _00778_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__12839__A _00392_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07644_ _05456_ VGND VGND VPWR VPWR _06417_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_95_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_832 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07575_ _05621_ _05544_ VGND VGND VPWR VPWR _05676_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_48_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09314_ _01332_ _01335_ VGND VGND VPWR VPWR _01457_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10078__B _02293_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09245_ _05566_ _00373_ _01089_ _01088_ VGND VGND VPWR VPWR _01382_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_63_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08670__A2 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_334 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_291 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09176_ _01245_ _01305_ VGND VGND VPWR VPWR _01307_ sky130_fd_sc_hd__nor2_4
XFILLER_0_133_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12293__B _01664_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12754__A1 _01504_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08127_ _00046_ _00073_ _00072_ VGND VGND VPWR VPWR _00171_ sky130_fd_sc_hd__a21bo_1
XANTENNA__12754__B2 _01507_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08058_ _00628_ _00650_ _00101_ _06733_ VGND VGND VPWR VPWR _00102_ sky130_fd_sc_hd__and4_1
XFILLER_0_101_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10822__A _03587_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput69 net69 VGND VGND VPWR VPWR prod[13] sky130_fd_sc_hd__clkbuf_4
X_10020_ _02229_ _02230_ VGND VGND VPWR VPWR _02231_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_399 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11971_ _04371_ _04372_ VGND VGND VPWR VPWR _04373_ sky130_fd_sc_hd__and2_1
X_13710_ _02759_ _05887_ _06267_ VGND VGND VPWR VPWR _06268_ sky130_fd_sc_hd__and3_1
X_10922_ _03215_ _03219_ VGND VGND VPWR VPWR _03220_ sky130_fd_sc_hd__nor2_1
XANTENNA__08894__C1 _00298_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13641_ _05975_ _05976_ VGND VGND VPWR VPWR _06192_ sky130_fd_sc_hd__or2_1
X_10853_ _03142_ _03143_ VGND VGND VPWR VPWR _03144_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13572_ _06114_ _06115_ VGND VGND VPWR VPWR _06116_ sky130_fd_sc_hd__nor2_2
XFILLER_0_67_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10784_ _03064_ _03067_ VGND VGND VPWR VPWR _03068_ sky130_fd_sc_hd__nand2_1
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12523_ _04944_ _04979_ VGND VGND VPWR VPWR _04980_ sky130_fd_sc_hd__and2b_1
XANTENNA__11796__A2 _02459_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_846 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12454_ _04883_ _04885_ VGND VGND VPWR VPWR _04904_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11548__A2 _02119_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11405_ _02119_ VGND VGND VPWR VPWR _03750_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_105_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12385_ _00778_ _00571_ _00734_ _00782_ VGND VGND VPWR VPWR _04828_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07728__D net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14124_ _06679_ _06682_ _06677_ VGND VGND VPWR VPWR _06721_ sky130_fd_sc_hd__o21ai_1
X_11336_ _03626_ _03667_ _03674_ VGND VGND VPWR VPWR _03675_ sky130_fd_sc_hd__and3_1
XFILLER_0_105_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14055_ _06613_ _06617_ _06620_ _06646_ VGND VGND VPWR VPWR _06647_ sky130_fd_sc_hd__o211a_1
X_11267_ _03531_ _03530_ _03518_ VGND VGND VPWR VPWR _03600_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_120_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13006_ _04602_ _04606_ _03578_ VGND VGND VPWR VPWR _05512_ sky130_fd_sc_hd__a21o_1
X_10218_ _05731_ _01177_ _01246_ _01000_ VGND VGND VPWR VPWR _02448_ sky130_fd_sc_hd__a22o_1
XANTENNA__11547__B _06966_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11198_ _03419_ _03438_ _03440_ VGND VGND VPWR VPWR _03524_ sky130_fd_sc_hd__a21oi_2
X_10149_ _02230_ _02371_ VGND VGND VPWR VPWR _02372_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13908_ _06433_ _06482_ _06485_ VGND VGND VPWR VPWR _06486_ sky130_fd_sc_hd__o21a_1
XANTENNA__13481__C _01958_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13839_ _06382_ _06385_ VGND VGND VPWR VPWR _06410_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_147_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_539 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07360_ _03290_ _03301_ VGND VGND VPWR VPWR _03312_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_742 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07291_ _02532_ _02543_ VGND VGND VPWR VPWR _02554_ sky130_fd_sc_hd__and2b_1
XFILLER_0_45_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08591__B _00523_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09030_ _01005_ _01146_ VGND VGND VPWR VPWR _01147_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07919__C net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_294 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12841__B _02168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09932_ _02133_ VGND VGND VPWR VPWR _02134_ sky130_fd_sc_hd__buf_2
XFILLER_0_111_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09863_ _02026_ _02057_ VGND VGND VPWR VPWR _02058_ sky130_fd_sc_hd__nand2_1
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08814_ _00738_ _00909_ VGND VGND VPWR VPWR _00910_ sky130_fd_sc_hd__nor2_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09794_ _06417_ _00574_ _01600_ _06439_ VGND VGND VPWR VPWR _01983_ sky130_fd_sc_hd__a22o_1
X_08745_ _00833_ _00834_ VGND VGND VPWR VPWR _00835_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09668__A1 _00654_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10278__A2 net53 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08676_ _00591_ _00757_ VGND VGND VPWR VPWR _00760_ sky130_fd_sc_hd__and2_1
XANTENNA__13391__C _03681_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07627_ _06197_ _06219_ _01996_ _03268_ VGND VGND VPWR VPWR _06230_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_95_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10089__A _02158_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_854 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07558_ _05478_ _01383_ VGND VGND VPWR VPWR _05489_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09597__B net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07489_ _04642_ _04708_ _04719_ VGND VGND VPWR VPWR _04730_ sky130_fd_sc_hd__or3_4
XFILLER_0_63_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09228_ _04048_ _01363_ VGND VGND VPWR VPWR _01364_ sky130_fd_sc_hd__and2_1
XANTENNA__07398__A _03718_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09159_ _00575_ VGND VGND VPWR VPWR _01288_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_133_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10738__B1 _02720_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12170_ _04548_ _04550_ VGND VGND VPWR VPWR _04592_ sky130_fd_sc_hd__nor2_1
XANTENNA__13847__B _03783_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11121_ _03396_ _03401_ _03388_ VGND VGND VPWR VPWR _03439_ sky130_fd_sc_hd__o21a_1
XFILLER_0_7_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_686 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11052_ _03351_ _03361_ _03362_ VGND VGND VPWR VPWR _03363_ sky130_fd_sc_hd__o21a_1
XANTENNA__10271__B _02308_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10003_ _05181_ _04037_ _01876_ _01874_ VGND VGND VPWR VPWR _02212_ sky130_fd_sc_hd__a31o_1
XANTENNA__08957__A _02467_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13582__B _03785_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11954_ _04282_ _04102_ _04283_ VGND VGND VPWR VPWR _04354_ sky130_fd_sc_hd__or3_2
X_10905_ _03082_ _03200_ VGND VGND VPWR VPWR _03201_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11885_ _04272_ _04277_ VGND VGND VPWR VPWR _04278_ sky130_fd_sc_hd__nor2_1
XANTENNA_output108_A net108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13624_ _06170_ _06172_ VGND VGND VPWR VPWR _06173_ sky130_fd_sc_hd__nand2_1
X_10836_ _01339_ _01933_ _02513_ VGND VGND VPWR VPWR _03126_ sky130_fd_sc_hd__and3_1
XANTENNA__09788__A _02456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08692__A net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11769__A2 _01564_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13555_ _06095_ _06096_ VGND VGND VPWR VPWR _06097_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10767_ _03016_ _03045_ _03049_ VGND VGND VPWR VPWR _03050_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_109_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12506_ _04959_ _04960_ VGND VGND VPWR VPWR _04962_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_42_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13486_ _06019_ _06020_ VGND VGND VPWR VPWR _06022_ sky130_fd_sc_hd__and2b_1
XFILLER_0_124_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10698_ _02965_ _02970_ _02972_ VGND VGND VPWR VPWR _02974_ sky130_fd_sc_hd__nand3_1
XFILLER_0_89_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_14 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07101__A net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12437_ _04883_ _04885_ VGND VGND VPWR VPWR _04886_ sky130_fd_sc_hd__or2_1
XFILLER_0_140_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12368_ _04793_ _04790_ VGND VGND VPWR VPWR _04810_ sky130_fd_sc_hd__xnor2_1
X_14107_ _06078_ _02742_ _06702_ VGND VGND VPWR VPWR _06703_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_1_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11319_ _03648_ _03656_ VGND VGND VPWR VPWR _03657_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07755__B _00508_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13476__C _01956_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12299_ _02188_ _02427_ VGND VGND VPWR VPWR _04734_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14038_ _06579_ _06618_ _06573_ VGND VGND VPWR VPWR _06629_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_38_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08570__A1 _06965_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08570__B2 _00263_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08530_ _00453_ _00460_ _00456_ _02467_ _00380_ VGND VGND VPWR VPWR _00600_ sky130_fd_sc_hd__a32o_1
XANTENNA__07490__B _04367_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08461_ _00466_ _00524_ VGND VGND VPWR VPWR _00525_ sky130_fd_sc_hd__xor2_1
XFILLER_0_77_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11443__D _02459_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07412_ _03861_ _03872_ VGND VGND VPWR VPWR _03883_ sky130_fd_sc_hd__and2b_1
XFILLER_0_9_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12406__B1 _00571_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08392_ _00447_ _00448_ VGND VGND VPWR VPWR _00449_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_147_347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07343_ _02576_ _02521_ VGND VGND VPWR VPWR _03125_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10637__A _01472_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09210__B _01343_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07274_ _02072_ _02083_ VGND VGND VPWR VPWR _02368_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08107__A _05181_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09013_ _01122_ _01127_ VGND VGND VPWR VPWR _01128_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_116_778 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08389__A1 _00880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__08389__B2 _04169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11393__B1 _01249_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11468__A _00497_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07665__B _06637_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09915_ _02138_ _01960_ _01968_ _01967_ VGND VGND VPWR VPWR _02115_ sky130_fd_sc_hd__a31o_1
XANTENNA__10091__B _02305_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09846_ _01951_ _02039_ VGND VGND VPWR VPWR _02041_ sky130_fd_sc_hd__xnor2_4
XANTENNA__11696__A1 _06873_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11696__B2 _06875_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07681__A net1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09777_ _01295_ _01246_ VGND VGND VPWR VPWR _01965_ sky130_fd_sc_hd__nand2_1
XANTENNA__12299__A _02188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08728_ _00643_ _00646_ VGND VGND VPWR VPWR _00817_ sky130_fd_sc_hd__and2_1
XTAP_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08659_ _03938_ VGND VGND VPWR VPWR _00741_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11353__D _03687_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11931__A _00113_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10671__A2 _02849_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11670_ _07010_ net38 _03718_ net10 VGND VGND VPWR VPWR _04042_ sky130_fd_sc_hd__and4_1
XANTENNA__10232__A1_N _00322_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10621_ _02876_ _02888_ VGND VGND VPWR VPWR _02889_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10547__A _00819_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13340_ _05326_ _05331_ VGND VGND VPWR VPWR _05862_ sky130_fd_sc_hd__and2_1
XFILLER_0_134_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07824__B1 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10552_ _02805_ _02812_ VGND VGND VPWR VPWR _02813_ sky130_fd_sc_hd__xor2_1
XANTENNA__10423__A2 net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11620__A1 _00544_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13271_ _05773_ _05776_ _05794_ VGND VGND VPWR VPWR _05795_ sky130_fd_sc_hd__a21o_1
XFILLER_0_122_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10483_ _02731_ VGND VGND VPWR VPWR _02737_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_122_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12222_ _04647_ _04648_ VGND VGND VPWR VPWR _04649_ sky130_fd_sc_hd__or2_1
XANTENNA__13577__B _02855_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12153_ _04570_ _04571_ _04572_ VGND VGND VPWR VPWR _04573_ sky130_fd_sc_hd__a21o_1
XFILLER_0_20_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11104_ _03412_ _03413_ VGND VGND VPWR VPWR _03420_ sky130_fd_sc_hd__or2_1
X_12084_ _04416_ _04419_ _04496_ VGND VGND VPWR VPWR _04497_ sky130_fd_sc_hd__o21a_1
X_11035_ _00298_ _01517_ _03343_ VGND VGND VPWR VPWR _03344_ sky130_fd_sc_hd__and3_1
XANTENNA__14201__B _00410_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12986_ _05485_ _05487_ _05488_ VGND VGND VPWR VPWR _05490_ sky130_fd_sc_hd__o21ai_4
X_11937_ _04333_ _04335_ VGND VGND VPWR VPWR _04336_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11868_ _04258_ _04259_ _00003_ _01600_ VGND VGND VPWR VPWR _04260_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_27_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10819_ _03105_ _03072_ _03101_ VGND VGND VPWR VPWR _03107_ sky130_fd_sc_hd__nor3_1
X_13607_ _01061_ _03785_ VGND VGND VPWR VPWR _06155_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_120 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11799_ _04182_ _04183_ VGND VGND VPWR VPWR _04184_ sky130_fd_sc_hd__nor2_1
X_13538_ _06074_ _06075_ _06077_ _06078_ VGND VGND VPWR VPWR _06079_ sky130_fd_sc_hd__and4_1
XFILLER_0_137_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13469_ _05994_ _06001_ VGND VGND VPWR VPWR _06003_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13364__A1 _01289_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13364__B2 _02008_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12391__B _01601_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09981__A _02187_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07961_ _02259_ _00004_ _07004_ _02171_ VGND VGND VPWR VPWR _00005_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_10_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09700_ _01870_ _01871_ _01879_ VGND VGND VPWR VPWR _01880_ sky130_fd_sc_hd__o21a_1
X_07892_ _00541_ _03499_ _06941_ _06940_ VGND VGND VPWR VPWR _07021_ sky130_fd_sc_hd__a31o_1
XANTENNA__08543__A1 _01230_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07346__A2 _00880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08543__B2 _01284_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09631_ _01610_ _01612_ _01804_ VGND VGND VPWR VPWR _01805_ sky130_fd_sc_hd__a21bo_1
XANTENNA__07932__C net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10350__A1 _02496_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13419__A2 _01415_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09562_ _00543_ _00859_ _01728_ VGND VGND VPWR VPWR _01729_ sky130_fd_sc_hd__and3_1
XFILLER_0_78_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08513_ _01295_ _03894_ _03938_ _01405_ VGND VGND VPWR VPWR _00581_ sky130_fd_sc_hd__a22o_1
X_09493_ _01372_ net50 VGND VGND VPWR VPWR _01653_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08444_ _00304_ _00306_ _00504_ VGND VGND VPWR VPWR _00506_ sky130_fd_sc_hd__nor3_1
XFILLER_0_93_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08375_ _00418_ _00419_ _00428_ VGND VGND VPWR VPWR _00430_ sky130_fd_sc_hd__nand3_1
XFILLER_0_73_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07326_ _00464_ _00530_ _02916_ VGND VGND VPWR VPWR _02938_ sky130_fd_sc_hd__and3_1
XFILLER_0_60_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07257_ _02116_ _02138_ _00333_ _02171_ VGND VGND VPWR VPWR _02182_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_5_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07676__A _06733_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07188_ _01350_ _01361_ _01416_ VGND VGND VPWR VPWR _01427_ sky130_fd_sc_hd__and3_1
XANTENNA__09023__A2 _00298_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11669__A1 _06733_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11669__B2 _03696_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09829_ _02010_ _02011_ _02020_ VGND VGND VPWR VPWR _02022_ sky130_fd_sc_hd__or3_1
X_12840_ _05327_ _05328_ VGND VGND VPWR VPWR _05329_ sky130_fd_sc_hd__nor2_1
XTAP_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12771_ _04649_ _04699_ _05252_ VGND VGND VPWR VPWR _05253_ sky130_fd_sc_hd__a21oi_1
XTAP_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11722_ _04097_ _04093_ _04094_ VGND VGND VPWR VPWR _04099_ sky130_fd_sc_hd__nor3_1
XTAP_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_656 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11653_ _04021_ _04022_ VGND VGND VPWR VPWR _04023_ sky130_fd_sc_hd__nor2_1
XTAP_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_816 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10604_ _02851_ _02848_ VGND VGND VPWR VPWR _02870_ sky130_fd_sc_hd__and2b_1
XFILLER_0_36_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11584_ _03944_ _03946_ VGND VGND VPWR VPWR _03947_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09262__A2 _00460_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07289__C net61 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13323_ _05748_ _05646_ VGND VGND VPWR VPWR _05844_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10535_ _02768_ _02769_ VGND VGND VPWR VPWR _02794_ sky130_fd_sc_hd__or2_1
XFILLER_0_101_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13254_ _05505_ _05506_ VGND VGND VPWR VPWR _05778_ sky130_fd_sc_hd__or2b_2
X_10466_ _02713_ _02718_ VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__xor2_4
XFILLER_0_20_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12205_ _00374_ _00784_ _01953_ _02134_ VGND VGND VPWR VPWR _04630_ sky130_fd_sc_hd__and4_1
XFILLER_0_86_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13185_ _05206_ _05707_ VGND VGND VPWR VPWR _05708_ sky130_fd_sc_hd__and2_1
X_10397_ _02640_ _02643_ VGND VGND VPWR VPWR _02644_ sky130_fd_sc_hd__xnor2_2
XANTENNA__07736__D net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12136_ _04491_ _04553_ VGND VGND VPWR VPWR _04555_ sky130_fd_sc_hd__and2b_1
XANTENNA__09970__B1 _01413_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09009__C _00114_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10580__A1 _00143_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10580__B2 _04906_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12067_ _04465_ _04474_ _04478_ VGND VGND VPWR VPWR _04479_ sky130_fd_sc_hd__a21o_1
X_11018_ _03324_ _03325_ VGND VGND VPWR VPWR _03326_ sky130_fd_sc_hd__and2_1
XFILLER_0_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12969_ _05455_ _05470_ VGND VGND VPWR VPWR _05471_ sky130_fd_sc_hd__xnor2_4
XANTENNA__08864__B net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_143_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12386__B _00613_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13034__B1 _05541_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10187__A _03499_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10618__C _01060_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08160_ _00202_ _06998_ _00203_ VGND VGND VPWR VPWR _00204_ sky130_fd_sc_hd__and3_1
XFILLER_0_7_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07111_ _00563_ net28 _00573_ net44 VGND VGND VPWR VPWR _00584_ sky130_fd_sc_hd__and4_1
XFILLER_0_70_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08091_ _00038_ _00039_ VGND VGND VPWR VPWR _00135_ sky130_fd_sc_hd__nor2_1
XANTENNA__09695__B _04367_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11348__B1 _03687_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13010__B _05513_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_543 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12560__A2 _04714_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08993_ _01064_ _01105_ VGND VGND VPWR VPWR _01106_ sky130_fd_sc_hd__xor2_1
XANTENNA__11746__A _00543_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07944_ _06926_ _07071_ _07042_ VGND VGND VPWR VPWR _07073_ sky130_fd_sc_hd__nand3_1
XANTENNA__12890__A1_N _01954_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07875_ _06885_ VGND VGND VPWR VPWR _07004_ sky130_fd_sc_hd__buf_4
X_09614_ _01784_ _01785_ VGND VGND VPWR VPWR _01786_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09545_ _01498_ _01708_ VGND VGND VPWR VPWR _01710_ sky130_fd_sc_hd__nor2_1
XANTENNA__12577__A _00389_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09476_ _01633_ _01634_ VGND VGND VPWR VPWR _01636_ sky130_fd_sc_hd__and2_4
XFILLER_0_78_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08427_ _00255_ _00266_ _00282_ VGND VGND VPWR VPWR _00488_ sky130_fd_sc_hd__o21a_1
XFILLER_0_19_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08358_ _04334_ _00348_ VGND VGND VPWR VPWR _00412_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07309_ _02675_ _02740_ VGND VGND VPWR VPWR _02751_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_144_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08289_ _00497_ _00151_ VGND VGND VPWR VPWR _00337_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10320_ _02361_ _02557_ VGND VGND VPWR VPWR _02559_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_830 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10251_ _02388_ _02389_ _02482_ VGND VGND VPWR VPWR _02484_ sky130_fd_sc_hd__nand3_2
XFILLER_0_104_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12551__A2 _01188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10182_ _02060_ _02406_ VGND VGND VPWR VPWR _02408_ sky130_fd_sc_hd__nand2_1
XANTENNA__10560__A _00294_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12303__A2 _02187_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09126__A _01250_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13941_ _06226_ _06228_ VGND VGND VPWR VPWR _06522_ sky130_fd_sc_hd__and2_1
XFILLER_0_89_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13872_ _06392_ _06400_ VGND VGND VPWR VPWR _06446_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12823_ _05308_ _04725_ _05309_ VGND VGND VPWR VPWR _05310_ sky130_fd_sc_hd__a21oi_1
XANTENNA__13590__B _01250_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12754_ _01504_ _01179_ _01254_ _01507_ VGND VGND VPWR VPWR _05234_ sky130_fd_sc_hd__a22o_1
XTAP_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11705_ _02418_ _02629_ _04078_ _04079_ VGND VGND VPWR VPWR _04080_ sky130_fd_sc_hd__o31a_1
XTAP_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12685_ _05156_ _05145_ _05150_ VGND VGND VPWR VPWR _05158_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_37_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_760 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11636_ _03877_ _03888_ VGND VGND VPWR VPWR _04005_ sky130_fd_sc_hd__and2b_1
XFILLER_0_37_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07246__A1 _00442_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07246__B2 _02051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11567_ _03532_ _00497_ _01179_ _01254_ VGND VGND VPWR VPWR _03929_ sky130_fd_sc_hd__and4_1
XFILLER_0_123_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10250__B1 _02482_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13319__A1 _05792_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10518_ _01473_ _02722_ VGND VGND VPWR VPWR _02776_ sky130_fd_sc_hd__nand2_1
X_13306_ _05667_ _05677_ VGND VGND VPWR VPWR _05828_ sky130_fd_sc_hd__nor2_1
XFILLER_0_123_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11498_ _03849_ _03852_ VGND VGND VPWR VPWR _03853_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13237_ _02491_ _02713_ _05575_ _05579_ VGND VGND VPWR VPWR _05763_ sky130_fd_sc_hd__and4_1
XFILLER_0_21_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10449_ _02699_ _02700_ VGND VGND VPWR VPWR _02701_ sky130_fd_sc_hd__or2_2
XFILLER_0_122_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13168_ _05683_ _05689_ VGND VGND VPWR VPWR _05690_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12119_ _04534_ _04535_ VGND VGND VPWR VPWR _04536_ sky130_fd_sc_hd__xor2_4
X_13099_ _05613_ VGND VGND VPWR VPWR _05614_ sky130_fd_sc_hd__inv_2
XANTENNA__13484__C _01957_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09171__A1 _03554_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07660_ _06560_ _06571_ VGND VGND VPWR VPWR _06593_ sky130_fd_sc_hd__and2_1
XANTENNA__09171__B2 _00519_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_830 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07591_ _05818_ _05827_ VGND VGND VPWR VPWR _05837_ sky130_fd_sc_hd__and2b_1
XFILLER_0_48_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09330_ _01471_ _01474_ VGND VGND VPWR VPWR _01475_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_62_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10629__B _02735_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09261_ _00608_ VGND VGND VPWR VPWR _01400_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_47_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13005__B _05494_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11451__D _02133_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08212_ _00118_ _00117_ VGND VGND VPWR VPWR _00256_ sky130_fd_sc_hd__and2b_1
XFILLER_0_16_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09192_ _01318_ _01323_ VGND VGND VPWR VPWR _01324_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09226__A2 _00376_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08143_ _06998_ _06999_ VGND VGND VPWR VPWR _00187_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07788__A2 _04367_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08074_ _00016_ _00018_ _00014_ VGND VGND VPWR VPWR _00118_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_70_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08115__A _01405_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08737__A1 _00258_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09934__B1 _02135_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10544__A1 _00819_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11476__A _03554_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10380__A _00486_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08976_ _00639_ net29 _04180_ _04191_ VGND VGND VPWR VPWR _01088_ sky130_fd_sc_hd__and4_1
X_07927_ _06905_ _06906_ VGND VGND VPWR VPWR _07056_ sky130_fd_sc_hd__nand2_1
XANTENNA__13691__A _02088_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07858_ _06898_ _06897_ _05412_ VGND VGND VPWR VPWR _06987_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08000__D _04939_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07789_ net59 _04455_ VGND VGND VPWR VPWR _06918_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09528_ _01690_ _01691_ VGND VGND VPWR VPWR _01692_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09459_ net64 _06820_ net8 net9 VGND VGND VPWR VPWR _01617_ sky130_fd_sc_hd__and4_1
XFILLER_0_66_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12470_ _02008_ _03414_ _01289_ _04714_ VGND VGND VPWR VPWR _04922_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_124_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11421_ _03765_ _03767_ VGND VGND VPWR VPWR _03768_ sky130_fd_sc_hd__and2b_1
XFILLER_0_123_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14140_ _06700_ _06710_ VGND VGND VPWR VPWR _06738_ sky130_fd_sc_hd__or2b_1
X_11352_ _01155_ _03680_ _03691_ VGND VGND VPWR VPWR _03692_ sky130_fd_sc_hd__and3_1
XFILLER_0_105_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10303_ _02180_ _02333_ _02539_ VGND VGND VPWR VPWR _02540_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_21_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14071_ _06077_ _04014_ _06662_ _06663_ VGND VGND VPWR VPWR _06664_ sky130_fd_sc_hd__o2bb2a_1
X_11283_ _03597_ _03601_ VGND VGND VPWR VPWR _03617_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13022_ _05510_ _05516_ VGND VGND VPWR VPWR _05529_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10234_ _02463_ _02464_ VGND VGND VPWR VPWR _02465_ sky130_fd_sc_hd__or2_1
X_10165_ _02387_ _02296_ _02298_ VGND VGND VPWR VPWR _02389_ sky130_fd_sc_hd__nand3_2
XANTENNA__13485__B1 _03690_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10096_ _00989_ net54 _02312_ _03576_ VGND VGND VPWR VPWR _02314_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13924_ _06499_ _06500_ _06502_ VGND VGND VPWR VPWR _06503_ sky130_fd_sc_hd__o21a_1
XANTENNA__07703__A2 net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13855_ _06424_ _06425_ VGND VGND VPWR VPWR _06427_ sky130_fd_sc_hd__xor2_1
XFILLER_0_85_800 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12806_ _05288_ _05054_ _05289_ _05290_ VGND VGND VPWR VPWR _05292_ sky130_fd_sc_hd__nand4_2
X_10998_ _03302_ _03269_ _03298_ VGND VGND VPWR VPWR _03304_ sky130_fd_sc_hd__nor3_1
X_13786_ _06349_ _05897_ _06350_ VGND VGND VPWR VPWR _06352_ sky130_fd_sc_hd__a21o_1
XFILLER_0_29_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07104__A _00497_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07467__A1 _00661_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12737_ _05171_ _05212_ _05215_ VGND VGND VPWR VPWR _05216_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_29_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12668_ _05132_ _05139_ VGND VGND VPWR VPWR _05140_ sky130_fd_sc_hd__or2b_1
XFILLER_0_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11619_ _03985_ _03932_ VGND VGND VPWR VPWR _03986_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_142_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12599_ _00914_ _01059_ _05062_ _05063_ VGND VGND VPWR VPWR _05064_ sky130_fd_sc_hd__a31o_1
XFILLER_0_25_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07196__D _01208_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07774__A _01470_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11296__A _00819_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08830_ _00924_ _00927_ VGND VGND VPWR VPWR _00928_ sky130_fd_sc_hd__xnor2_1
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08761_ _00851_ _00852_ VGND VGND VPWR VPWR _00853_ sky130_fd_sc_hd__nor2_2
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07712_ _06833_ _06839_ _06840_ VGND VGND VPWR VPWR _06841_ sky130_fd_sc_hd__or3_1
X_08692_ net43 VGND VGND VPWR VPWR _00777_ sky130_fd_sc_hd__buf_2
XANTENNA__12839__B _00742_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07643_ _06384_ _06395_ VGND VGND VPWR VPWR _06406_ sky130_fd_sc_hd__or2b_1
XANTENNA__13016__A _05501_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07574_ _05522_ _05533_ _05632_ _05643_ VGND VGND VPWR VPWR _05665_ sky130_fd_sc_hd__or4_4
XFILLER_0_76_844 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09313_ _01454_ _01455_ VGND VGND VPWR VPWR _01456_ sky130_fd_sc_hd__nor2_1
XANTENNA__07458__A1 net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12855__A _01584_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09244_ _01085_ _01093_ VGND VGND VPWR VPWR _01381_ sky130_fd_sc_hd__and2b_1
XFILLER_0_8_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09175_ _01256_ _01304_ VGND VGND VPWR VPWR _01305_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_113_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12293__C _01601_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08126_ _00150_ _00168_ _00169_ _00166_ VGND VGND VPWR VPWR _00170_ sky130_fd_sc_hd__o22a_1
XFILLER_0_44_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12754__A2 _01179_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10765__A1 _01156_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08057_ net38 VGND VGND VPWR VPWR _00101_ sky130_fd_sc_hd__buf_2
XANTENNA__13686__A _02427_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12590__A _00915_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10822__B _00891_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08959_ _00971_ _00974_ _00957_ VGND VGND VPWR VPWR _01069_ sky130_fd_sc_hd__o21a_1
X_11970_ _04369_ _04370_ _04303_ VGND VGND VPWR VPWR _04372_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09404__A _01500_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10921_ _03216_ _03218_ VGND VGND VPWR VPWR _03219_ sky130_fd_sc_hd__and2b_1
XANTENNA__08894__B1 _00508_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13640_ _06172_ _06190_ VGND VGND VPWR VPWR _06191_ sky130_fd_sc_hd__xor2_1
XFILLER_0_39_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10852_ _03268_ _02158_ _02304_ _05577_ VGND VGND VPWR VPWR _03143_ sky130_fd_sc_hd__a22oi_1
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13571_ _06113_ _06083_ VGND VGND VPWR VPWR _06115_ sky130_fd_sc_hd__and2b_1
XFILLER_0_137_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10783_ _03065_ _03066_ VGND VGND VPWR VPWR _03067_ sky130_fd_sc_hd__nor2_1
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10453__B1 _02703_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12522_ _04954_ _04977_ _04978_ VGND VGND VPWR VPWR _04979_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_137_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12453_ _04900_ _04902_ VGND VGND VPWR VPWR _04903_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11404_ _00004_ _03748_ _03742_ _03741_ VGND VGND VPWR VPWR _03749_ sky130_fd_sc_hd__a31o_1
XFILLER_0_50_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12384_ _04778_ _04787_ _04826_ VGND VGND VPWR VPWR _04827_ sky130_fd_sc_hd__and3_1
XFILLER_0_62_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_446 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14123_ _06719_ VGND VGND VPWR VPWR _06720_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11335_ _03673_ VGND VGND VPWR VPWR _03674_ sky130_fd_sc_hd__inv_2
XFILLER_0_132_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11266_ _03531_ _03518_ _03530_ VGND VGND VPWR VPWR _03599_ sky130_fd_sc_hd__or3_1
X_14054_ _06628_ _06645_ VGND VGND VPWR VPWR _06646_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13005_ _05493_ _05494_ VGND VGND VPWR VPWR _05510_ sky130_fd_sc_hd__xor2_2
X_10217_ _02444_ _02446_ VGND VGND VPWR VPWR _02447_ sky130_fd_sc_hd__xnor2_2
X_11197_ _03519_ _03522_ VGND VGND VPWR VPWR _03523_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_94_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11547__C _02119_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10148_ _02367_ _02370_ VGND VGND VPWR VPWR _02371_ sky130_fd_sc_hd__nor2_1
X_10079_ _02282_ _02293_ VGND VGND VPWR VPWR _02295_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13907_ _06414_ _06484_ VGND VGND VPWR VPWR _06485_ sky130_fd_sc_hd__nor2_1
XANTENNA__07688__A1 _01120_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13481__D _03690_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13838_ _06401_ _06408_ _06405_ VGND VGND VPWR VPWR _06409_ sky130_fd_sc_hd__o21a_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10179__B _03894_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_77 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13769_ _06316_ _06319_ VGND VGND VPWR VPWR _06333_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07290_ net62 _00923_ net61 _00869_ VGND VGND VPWR VPWR _02543_ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09344__C_N _01486_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09931_ net22 VGND VGND VPWR VPWR _02133_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_68_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09862_ _00519_ _01188_ _02025_ VGND VGND VPWR VPWR _02057_ sky130_fd_sc_hd__a21o_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08813_ _00905_ _00908_ VGND VGND VPWR VPWR _00909_ sky130_fd_sc_hd__xnor2_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09793_ _01774_ _01778_ _01775_ VGND VGND VPWR VPWR _01982_ sky130_fd_sc_hd__o21ba_1
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08744_ _00824_ _00832_ VGND VGND VPWR VPWR _00834_ sky130_fd_sc_hd__or2_1
XANTENNA__09668__A2 _00859_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08675_ _00591_ _00757_ VGND VGND VPWR VPWR _00758_ sky130_fd_sc_hd__nor2_1
XANTENNA__13391__D _02673_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07626_ _05445_ _00650_ _06208_ VGND VGND VPWR VPWR _06219_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_67_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08628__B1 _00547_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07557_ _05467_ VGND VGND VPWR VPWR _05478_ sky130_fd_sc_hd__buf_4
XFILLER_0_48_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_140 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07488_ _04411_ _04477_ VGND VGND VPWR VPWR _04719_ sky130_fd_sc_hd__xor2_1
XFILLER_0_90_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09227_ _00355_ _02960_ _04015_ VGND VGND VPWR VPWR _01363_ sky130_fd_sc_hd__and3_1
XFILLER_0_51_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09158_ _01285_ _01286_ VGND VGND VPWR VPWR _01287_ sky130_fd_sc_hd__nand2_1
XANTENNA__09894__A _06626_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10738__A1 _03015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10738__B2 _00399_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08109_ _06417_ _00151_ _00152_ VGND VGND VPWR VPWR _00153_ sky130_fd_sc_hd__and3_1
XFILLER_0_121_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09089_ _01209_ _01210_ _01744_ _01211_ VGND VGND VPWR VPWR _01212_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_114_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11120_ _03430_ _03434_ _03436_ _03437_ VGND VGND VPWR VPWR _03438_ sky130_fd_sc_hd__a31o_2
XFILLER_0_101_120 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11051_ _03342_ _03344_ VGND VGND VPWR VPWR _03362_ sky130_fd_sc_hd__xor2_1
XFILLER_0_102_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10002_ _01872_ _01878_ VGND VGND VPWR VPWR _02211_ sky130_fd_sc_hd__nand2_1
XANTENNA__08957__B _01066_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13582__C _02858_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09134__A _03938_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11953_ _04351_ _04352_ VGND VGND VPWR VPWR _04353_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10904_ _03079_ _03080_ VGND VGND VPWR VPWR _03200_ sky130_fd_sc_hd__or2_1
X_11884_ _04274_ _04276_ VGND VGND VPWR VPWR _04277_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_129_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13623_ _06031_ _06171_ VGND VGND VPWR VPWR _06172_ sky130_fd_sc_hd__or2_1
X_10835_ _03119_ _03122_ _03123_ VGND VGND VPWR VPWR _03124_ sky130_fd_sc_hd__and3_1
XFILLER_0_104_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09788__B _01180_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12495__A _04037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07589__A _05445_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13554_ _06092_ _06068_ _06094_ VGND VGND VPWR VPWR _06096_ sky130_fd_sc_hd__o21a_1
XFILLER_0_13_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10766_ _03046_ _03047_ VGND VGND VPWR VPWR _03049_ sky130_fd_sc_hd__nand2_1
XFILLER_0_137_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12505_ _04037_ _03773_ VGND VGND VPWR VPWR _04960_ sky130_fd_sc_hd__nand2_1
XFILLER_0_124_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07842__A1 _06967_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13485_ _06018_ _01957_ _03690_ _06009_ VGND VGND VPWR VPWR _06020_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10697_ _02965_ _02970_ _02972_ VGND VGND VPWR VPWR _02973_ sky130_fd_sc_hd__a21o_1
XFILLER_0_23_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12436_ _04837_ _04872_ VGND VGND VPWR VPWR _04885_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_112_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12367_ _04801_ _04806_ _04808_ VGND VGND VPWR VPWR _04809_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_22_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14106_ _02743_ _04014_ VGND VGND VPWR VPWR _06702_ sky130_fd_sc_hd__nand2_1
XANTENNA_output82_A net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09309__A _00843_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11318_ _03649_ _03646_ VGND VGND VPWR VPWR _03656_ sky130_fd_sc_hd__or2b_1
X_12298_ _04728_ _04732_ VGND VGND VPWR VPWR _04733_ sky130_fd_sc_hd__and2_1
XANTENNA__13476__D _03687_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08213__A _00113_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09347__A1 _02960_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09347__B2 _00355_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11249_ _03566_ _03579_ VGND VGND VPWR VPWR _03580_ sky130_fd_sc_hd__xor2_1
X_14037_ _06623_ _06627_ VGND VGND VPWR VPWR _06628_ sky130_fd_sc_hd__or2b_1
XFILLER_0_129_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__07358__B1 _02719_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12351__B1 _01369_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__08570__A2 _00293_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07771__B _00573_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12654__A1 _00390_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08460_ _00493_ _00523_ VGND VGND VPWR VPWR _00524_ sky130_fd_sc_hd__xor2_2
XFILLER_0_58_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07411_ _03850_ _03685_ _03718_ _01306_ VGND VGND VPWR VPWR _03872_ sky130_fd_sc_hd__a22o_1
XFILLER_0_147_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08391_ _04268_ _04026_ VGND VGND VPWR VPWR _00448_ sky130_fd_sc_hd__nand2_1
XANTENNA__12406__A1 _00782_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12406__B2 _00373_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07342_ _03081_ _03103_ VGND VGND VPWR VPWR _03114_ sky130_fd_sc_hd__and2_1
XFILLER_0_57_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10637__B _02856_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_143_510 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07273_ _02270_ _02324_ _02346_ VGND VGND VPWR VPWR _02357_ sky130_fd_sc_hd__o21a_1
XFILLER_0_73_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09012_ _01125_ _01126_ VGND VGND VPWR VPWR _01127_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11393__A1 _00113_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11393__B2 _00114_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11468__B _02673_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09914_ _01964_ _01970_ VGND VGND VPWR VPWR _02114_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07962__A _02259_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09845_ _02036_ _02037_ _02038_ VGND VGND VPWR VPWR _02039_ sky130_fd_sc_hd__or3_4
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11696__A2 _01272_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07681__B net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09776_ _01178_ _01808_ _01811_ _01812_ VGND VGND VPWR VPWR _01964_ sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__12299__B _02427_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08727_ _00813_ _00815_ VGND VGND VPWR VPWR _00816_ sky130_fd_sc_hd__nand2_1
XTAP_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08658_ _00738_ _00739_ VGND VGND VPWR VPWR _00740_ sky130_fd_sc_hd__and2_2
XFILLER_0_96_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07609_ _05808_ _06021_ VGND VGND VPWR VPWR _06032_ sky130_fd_sc_hd__nand2_2
XFILLER_0_49_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11931__B _00114_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10828__A _01383_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08589_ _00634_ _00663_ VGND VGND VPWR VPWR _00665_ sky130_fd_sc_hd__and2_1
X_10620_ _02873_ _02875_ VGND VGND VPWR VPWR _02888_ sky130_fd_sc_hd__or2_1
XFILLER_0_76_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10959__A1 _00859_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10547__B _00818_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07202__A _01230_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07824__A1 _00420_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10551_ _02810_ _02811_ VGND VGND VPWR VPWR _02812_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11620__A2 _01182_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07824__B2 net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_705 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13270_ _05779_ _05793_ VGND VGND VPWR VPWR _05794_ sky130_fd_sc_hd__nand2_1
X_10482_ _02735_ VGND VGND VPWR VPWR _02736_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_134_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12221_ _04645_ _04646_ VGND VGND VPWR VPWR _04648_ sky130_fd_sc_hd__and2_1
XANTENNA__13577__C _03785_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12581__B1 _02304_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12152_ _02694_ _02698_ VGND VGND VPWR VPWR _04572_ sky130_fd_sc_hd__nand2_1
XANTENNA__09129__A _02138_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11103_ _03404_ _03418_ VGND VGND VPWR VPWR _03419_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_102_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12083_ _04494_ _04495_ VGND VGND VPWR VPWR _04496_ sky130_fd_sc_hd__nor2_1
XANTENNA__07872__A _00530_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11034_ _00143_ _01518_ VGND VGND VPWR VPWR _03343_ sky130_fd_sc_hd__nand2_1
XANTENNA__11394__A _02119_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output120_A net120 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12985_ _05476_ _05484_ VGND VGND VPWR VPWR _05488_ sky130_fd_sc_hd__or2_1
X_11936_ _00004_ _01585_ _04332_ VGND VGND VPWR VPWR _04335_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_129_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11867_ _00113_ _00415_ _00575_ _00258_ VGND VGND VPWR VPWR _04259_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_28_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13606_ _02856_ _06145_ _06144_ VGND VGND VPWR VPWR _06154_ sky130_fd_sc_hd__a21bo_1
X_10818_ _03072_ _03101_ _03105_ VGND VGND VPWR VPWR _03106_ sky130_fd_sc_hd__o21a_1
XFILLER_0_144_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11798_ _04179_ _04181_ _04173_ _04175_ VGND VGND VPWR VPWR _04183_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_28_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13537_ _03690_ VGND VGND VPWR VPWR _06078_ sky130_fd_sc_hd__buf_2
XFILLER_0_15_519 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10749_ _03025_ _03028_ VGND VGND VPWR VPWR _03030_ sky130_fd_sc_hd__nor2_1
XFILLER_0_131_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13468_ _05994_ _06001_ VGND VGND VPWR VPWR _06002_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12419_ _04864_ _04865_ VGND VGND VPWR VPWR _04866_ sky130_fd_sc_hd__and2b_1
XANTENNA__13364__A2 _02759_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10473__A _02725_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13399_ _05925_ _05926_ VGND VGND VPWR VPWR _05927_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07960_ _00003_ VGND VGND VPWR VPWR _00004_ sky130_fd_sc_hd__clkbuf_4
X_07891_ _06944_ _06947_ _07019_ VGND VGND VPWR VPWR _07020_ sky130_fd_sc_hd__a21o_1
XFILLER_0_65_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08543__A2 _00612_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09630_ _01608_ _01609_ VGND VGND VPWR VPWR _01804_ sky130_fd_sc_hd__or2b_1
XANTENNA__10350__A2 _02498_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07932__D net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09415__A2_N _01564_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09561_ _00543_ _01472_ _01469_ _01468_ _07040_ VGND VGND VPWR VPWR _01728_ sky130_fd_sc_hd__a32o_1
X_08512_ _00421_ _00427_ VGND VGND VPWR VPWR _00580_ sky130_fd_sc_hd__nand2_1
X_09492_ _01650_ _01651_ VGND VGND VPWR VPWR _01652_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08443_ _00304_ _00306_ _00504_ VGND VGND VPWR VPWR _00505_ sky130_fd_sc_hd__o21a_1
XFILLER_0_58_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08374_ _00418_ _00419_ _00428_ VGND VGND VPWR VPWR _00429_ sky130_fd_sc_hd__a21o_1
XFILLER_0_45_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07325_ _00464_ _00530_ _02916_ VGND VGND VPWR VPWR _02927_ sky130_fd_sc_hd__a21o_1
XFILLER_0_61_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07256_ _02160_ VGND VGND VPWR VPWR _02171_ sky130_fd_sc_hd__buf_4
XANTENNA__09008__B1 _00114_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07187_ _01383_ _01405_ VGND VGND VPWR VPWR _01416_ sky130_fd_sc_hd__nand2_1
XFILLER_0_131_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07692__A _06820_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11669__A2 _03773_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09828_ _02010_ _02011_ _02020_ VGND VGND VPWR VPWR _02021_ sky130_fd_sc_hd__o21a_1
X_09759_ _01942_ _01944_ VGND VGND VPWR VPWR _01945_ sky130_fd_sc_hd__xor2_1
XTAP_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12770_ _04649_ _04699_ _04638_ VGND VGND VPWR VPWR _05252_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_96_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ _04093_ _04094_ _04097_ VGND VGND VPWR VPWR _04098_ sky130_fd_sc_hd__o21a_1
XTAP_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10558__A _00293_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11652_ _04020_ _03844_ _04012_ VGND VGND VPWR VPWR _04022_ sky130_fd_sc_hd__and3_1
XTAP_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10603_ _02866_ _02868_ VGND VGND VPWR VPWR _02869_ sky130_fd_sc_hd__or2_1
XFILLER_0_92_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11583_ _03832_ _03945_ VGND VGND VPWR VPWR _03946_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_828 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07289__D _00869_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13322_ _05795_ _05798_ _05815_ _05842_ VGND VGND VPWR VPWR _05843_ sky130_fd_sc_hd__a211o_1
X_10534_ _02792_ VGND VGND VPWR VPWR _02793_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10465_ _01649_ _02275_ _02714_ _02717_ VGND VGND VPWR VPWR _02718_ sky130_fd_sc_hd__a31o_1
X_13253_ _05524_ net130 VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__xor2_4
XFILLER_0_122_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12204_ _04601_ _04628_ VGND VGND VPWR VPWR _04629_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13184_ _05202_ _05205_ VGND VGND VPWR VPWR _05707_ sky130_fd_sc_hd__nand2_1
X_10396_ _02082_ _02422_ _02641_ VGND VGND VPWR VPWR _02643_ sky130_fd_sc_hd__a21o_1
XFILLER_0_103_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12135_ _04537_ _04552_ VGND VGND VPWR VPWR _04553_ sky130_fd_sc_hd__nor2_1
XANTENNA__09970__A1 _02171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09970__B2 _02259_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08698__A _00783_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09009__D _00094_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10580__A2 _02306_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12066_ _04475_ _04476_ VGND VGND VPWR VPWR _04478_ sky130_fd_sc_hd__and2_1
X_11017_ _03316_ _03319_ VGND VGND VPWR VPWR _03325_ sky130_fd_sc_hd__xor2_1
XANTENNA__08210__B _00175_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07107__A net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_360 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12968_ _05457_ _05469_ VGND VGND VPWR VPWR _05470_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_59_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10096__A1 _00989_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11919_ _04305_ _04315_ VGND VGND VPWR VPWR _04316_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10096__B2 _03576_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10468__A _02720_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12899_ _05230_ _05393_ VGND VGND VPWR VPWR _05394_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_600 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_216 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12386__C _00571_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10187__B _06821_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09789__A1 _02456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10618__D _01413_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_772 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07110_ net55 VGND VGND VPWR VPWR _00573_ sky130_fd_sc_hd__buf_6
X_08090_ _00132_ _00133_ VGND VGND VPWR VPWR _00134_ sky130_fd_sc_hd__xnor2_2
XANTENNA__07777__A net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13601__A2_N _03785_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11348__A1 _02249_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11348__B2 _01312_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08992_ _01067_ _01104_ VGND VGND VPWR VPWR _01105_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_76_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07943_ _06926_ _07042_ _07071_ VGND VGND VPWR VPWR _07072_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11746__B _01188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08401__A _00458_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07874_ _06976_ _06979_ _07002_ VGND VGND VPWR VPWR _07003_ sky130_fd_sc_hd__a21o_1
XANTENNA__07724__B1 _00508_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09613_ _01782_ _01783_ _01779_ VGND VGND VPWR VPWR _01785_ sky130_fd_sc_hd__o21a_1
XFILLER_0_97_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11762__A _00138_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09544_ _01498_ _01708_ VGND VGND VPWR VPWR _01709_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12577__B _00393_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09232__A net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09475_ _01631_ _01632_ _01428_ _01431_ VGND VGND VPWR VPWR _01634_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_93_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08426_ _00484_ _00485_ VGND VGND VPWR VPWR _00487_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08357_ _00372_ _00411_ VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__xor2_2
XFILLER_0_74_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire129 net113 VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__buf_4
XFILLER_0_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07308_ _02708_ _02729_ VGND VGND VPWR VPWR _02740_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_116_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08288_ _00497_ _00094_ _00092_ _00091_ VGND VGND VPWR VPWR _00336_ sky130_fd_sc_hd__a31o_1
XFILLER_0_144_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07239_ _01886_ _01974_ VGND VGND VPWR VPWR _01985_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10250_ _02388_ _02389_ _02482_ VGND VGND VPWR VPWR _02483_ sky130_fd_sc_hd__a21o_1
XFILLER_0_30_842 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10181_ _02060_ _02406_ VGND VGND VPWR VPWR _02407_ sky130_fd_sc_hd__or2_2
XFILLER_0_100_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10560__B _01934_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13940_ _06509_ _06520_ VGND VGND VPWR VPWR _06521_ sky130_fd_sc_hd__xnor2_4
X_13871_ _06442_ _06444_ VGND VGND VPWR VPWR _06445_ sky130_fd_sc_hd__nand2_1
XANTENNA__11466__A2_N _03681_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12822_ _05039_ _05130_ VGND VGND VPWR VPWR _05309_ sky130_fd_sc_hd__nor2_1
XANTENNA__13590__C _02856_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09468__B1 _01626_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12753_ _01507_ _01504_ _01248_ VGND VGND VPWR VPWR _05233_ sky130_fd_sc_hd__and3_1
XANTENNA__10288__A _00628_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11704_ _04076_ _02627_ _04077_ VGND VGND VPWR VPWR _04079_ sky130_fd_sc_hd__a21o_1
XTAP_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12684_ _05156_ _05145_ _05150_ VGND VGND VPWR VPWR _05157_ sky130_fd_sc_hd__or3_1
XFILLER_0_139_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11635_ _03891_ _03954_ _04002_ VGND VGND VPWR VPWR _04003_ sky130_fd_sc_hd__o21bai_4
XFILLER_0_65_772 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_660 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07246__A2 _02018_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11566_ _03925_ _03926_ VGND VGND VPWR VPWR _03928_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_13_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13319__A2 _05807_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13305_ _05678_ _05694_ VGND VGND VPWR VPWR _05826_ sky130_fd_sc_hd__and2_1
XFILLER_0_107_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10517_ _02752_ _02750_ VGND VGND VPWR VPWR _02775_ sky130_fd_sc_hd__and2b_1
XFILLER_0_80_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11497_ _03840_ _03851_ VGND VGND VPWR VPWR _03852_ sky130_fd_sc_hd__and2_1
X_13236_ _05760_ VGND VGND VPWR VPWR _05762_ sky130_fd_sc_hd__inv_2
X_10448_ _02476_ _02480_ VGND VGND VPWR VPWR _02700_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13167_ _05685_ _05688_ VGND VGND VPWR VPWR _05689_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10379_ _00475_ _00734_ _02411_ _02414_ VGND VGND VPWR VPWR _02624_ sky130_fd_sc_hd__a31o_1
XFILLER_0_20_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12118_ _04451_ _04450_ VGND VGND VPWR VPWR _04535_ sky130_fd_sc_hd__and2b_2
X_13098_ _04025_ _04546_ VGND VGND VPWR VPWR _05613_ sky130_fd_sc_hd__or2_1
XANTENNA__13484__D _03690_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12049_ _04134_ _04137_ _04139_ VGND VGND VPWR VPWR _04459_ sky130_fd_sc_hd__and3_1
XFILLER_0_137_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09171__A2 _00391_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07590_ _05456_ _02105_ _00650_ _05467_ VGND VGND VPWR VPWR _05827_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_842 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10198__A _02088_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09260_ _02116_ _02160_ _00605_ VGND VGND VPWR VPWR _01399_ sky130_fd_sc_hd__and3_1
XFILLER_0_8_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08211_ _00119_ _00126_ VGND VGND VPWR VPWR _00255_ sky130_fd_sc_hd__nand2_1
XFILLER_0_118_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09191_ _01319_ _01322_ VGND VGND VPWR VPWR _01323_ sky130_fd_sc_hd__xor2_1
XFILLER_0_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10926__A _02467_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08142_ _00184_ _00185_ VGND VGND VPWR VPWR _00186_ sky130_fd_sc_hd__and2_1
XFILLER_0_71_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08073_ _00111_ _00116_ VGND VGND VPWR VPWR _00117_ sky130_fd_sc_hd__xor2_1
XFILLER_0_125_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09934__A1 _02138_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09934__B2 _00333_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10544__A2 _02169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09227__A _00355_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11476__B _00508_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08975_ _05577_ _00373_ _00946_ _00944_ VGND VGND VPWR VPWR _01086_ sky130_fd_sc_hd__a31o_1
XANTENNA__10380__B _01211_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07926_ _06921_ _07054_ VGND VGND VPWR VPWR _07055_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13691__B _02720_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07857_ _06898_ _05412_ _06897_ VGND VGND VPWR VPWR _06986_ sky130_fd_sc_hd__or3_4
XANTENNA__07173__A1 _01230_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07788_ net59 _04367_ _05104_ _05093_ VGND VGND VPWR VPWR _06917_ sky130_fd_sc_hd__a31o_1
XFILLER_0_79_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09527_ _01688_ _01686_ VGND VGND VPWR VPWR _01691_ sky130_fd_sc_hd__and2b_1
XFILLER_0_38_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09458_ _01615_ VGND VGND VPWR VPWR _01616_ sky130_fd_sc_hd__inv_2
X_08409_ _00288_ _00467_ _00286_ VGND VGND VPWR VPWR _00468_ sky130_fd_sc_hd__a21o_1
XFILLER_0_47_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10480__A1 _02247_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10836__A _01339_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09389_ _01396_ _01402_ _01397_ VGND VGND VPWR VPWR _01540_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_62_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11420_ _03763_ _03766_ VGND VGND VPWR VPWR _03767_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11351_ _00544_ _03684_ _03688_ _03689_ _03690_ VGND VGND VPWR VPWR _03691_ sky130_fd_sc_hd__a32o_1
XFILLER_0_34_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10302_ _02301_ _02332_ VGND VGND VPWR VPWR _02539_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_691 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14070_ _06075_ _06078_ _02743_ _02742_ VGND VGND VPWR VPWR _06663_ sky130_fd_sc_hd__and4_1
XFILLER_0_21_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11282_ _03585_ _03588_ _03590_ _03612_ _03615_ VGND VGND VPWR VPWR _03616_ sky130_fd_sc_hd__a311oi_2
XFILLER_0_120_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13021_ _02049_ _05526_ _05527_ _02492_ VGND VGND VPWR VPWR _05528_ sky130_fd_sc_hd__o31ai_4
XANTENNA__11667__A _00004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10233_ _02462_ net24 _00322_ _02460_ VGND VGND VPWR VPWR _02464_ sky130_fd_sc_hd__and4b_1
XFILLER_0_120_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10571__A _00399_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10164_ _02296_ _02298_ _02387_ VGND VGND VPWR VPWR _02388_ sky130_fd_sc_hd__a21o_1
X_10095_ net56 VGND VGND VPWR VPWR _02312_ sky130_fd_sc_hd__buf_2
XANTENNA__08976__A _00639_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13923_ _06203_ _06229_ VGND VGND VPWR VPWR _06502_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_107_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13854_ _06424_ _06425_ VGND VGND VPWR VPWR _06426_ sky130_fd_sc_hd__nand2_1
X_12805_ _05111_ _05113_ VGND VGND VPWR VPWR _05290_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13106__B _05620_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13785_ _06346_ _06347_ VGND VGND VPWR VPWR _06350_ sky130_fd_sc_hd__xor2_1
X_10997_ _03269_ _03298_ _03302_ VGND VGND VPWR VPWR _03303_ sky130_fd_sc_hd__o21a_1
XFILLER_0_123_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12736_ _05152_ _05213_ VGND VGND VPWR VPWR _05215_ sky130_fd_sc_hd__xnor2_1
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08664__A1 _00157_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12667_ _05133_ _05134_ _05138_ VGND VGND VPWR VPWR _05139_ sky130_fd_sc_hd__o21ba_1
XANTENNA__14218__A _00464_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11618_ _03933_ _03924_ VGND VGND VPWR VPWR _03985_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12598_ _03707_ _03740_ _01411_ _02849_ VGND VGND VPWR VPWR _05063_ sky130_fd_sc_hd__and4_1
XFILLER_0_114_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07120__A _00628_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11549_ _03906_ _03907_ _03908_ VGND VGND VPWR VPWR _03909_ sky130_fd_sc_hd__and3_1
XFILLER_0_123_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_639 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13219_ _05660_ _05662_ VGND VGND VPWR VPWR _05746_ sky130_fd_sc_hd__and2b_1
XFILLER_0_110_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10481__A _02726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07774__B net6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14199_ _02357_ _02390_ VGND VGND VPWR VPWR _06792_ sky130_fd_sc_hd__nor2_1
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11296__B _00818_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08760_ _00676_ _00681_ _00850_ VGND VGND VPWR VPWR _00852_ sky130_fd_sc_hd__o21a_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07711_ _06809_ _06816_ VGND VGND VPWR VPWR _06840_ sky130_fd_sc_hd__xor2_1
X_08691_ _00611_ _00616_ VGND VGND VPWR VPWR _00776_ sky130_fd_sc_hd__nor2_1
XANTENNA__12839__C _02723_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07642_ _06362_ _06373_ VGND VGND VPWR VPWR _06395_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07573_ net151 _05533_ _05632_ _05643_ VGND VGND VPWR VPWR _05654_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_88_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09312_ _01449_ _01327_ _01453_ VGND VGND VPWR VPWR _01455_ sky130_fd_sc_hd__o21a_1
XFILLER_0_75_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_856 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07458__A2 net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12855__B _01412_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09510__A _06494_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09243_ _01378_ _01379_ VGND VGND VPWR VPWR _01380_ sky130_fd_sc_hd__nor2_1
XFILLER_0_63_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09174_ _01300_ _01303_ VGND VGND VPWR VPWR _01304_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08125_ _00069_ _00165_ _00150_ VGND VGND VPWR VPWR _00169_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12293__D _01505_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11962__A1 _03059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10765__A2 _02766_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08056_ _00098_ _00099_ VGND VGND VPWR VPWR _00100_ sky130_fd_sc_hd__or2_2
XFILLER_0_98_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13686__B _02426_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12590__B _00916_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10822__C net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08958_ _00971_ _00974_ VGND VGND VPWR VPWR _01068_ sky130_fd_sc_hd__and2_1
X_07909_ _06931_ _06929_ VGND VGND VPWR VPWR _07038_ sky130_fd_sc_hd__and2b_1
XANTENNA__12675__C1 _01958_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08889_ _06965_ _06966_ _04906_ _04928_ VGND VGND VPWR VPWR _00993_ sky130_fd_sc_hd__and4_1
XANTENNA__08343__B1 _00395_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10920_ _03080_ _03217_ VGND VGND VPWR VPWR _03218_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10851_ _02664_ _03268_ _01546_ _02156_ VGND VGND VPWR VPWR _03142_ sky130_fd_sc_hd__and4_1
XFILLER_0_67_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13570_ _06083_ _06113_ VGND VGND VPWR VPWR _06114_ sky130_fd_sc_hd__and2b_1
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10782_ _06637_ _02726_ _02730_ _06937_ VGND VGND VPWR VPWR _03066_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_93_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12521_ _04947_ _04951_ _04953_ VGND VGND VPWR VPWR _04978_ sky130_fd_sc_hd__nand3_1
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12452_ _04901_ _04870_ VGND VGND VPWR VPWR _04902_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_136_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11403_ _03744_ VGND VGND VPWR VPWR _03748_ sky130_fd_sc_hd__clkbuf_4
X_12383_ _04798_ _04824_ _04825_ VGND VGND VPWR VPWR _04826_ sky130_fd_sc_hd__o21ai_1
X_14122_ _06716_ _06718_ VGND VGND VPWR VPWR _06719_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07875__A _06885_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11334_ _03668_ _03672_ VGND VGND VPWR VPWR _03673_ sky130_fd_sc_hd__or2_1
XFILLER_0_132_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_458 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14053_ _06632_ _06644_ VGND VGND VPWR VPWR _06645_ sky130_fd_sc_hd__or2_2
X_11265_ _03593_ _03595_ _03596_ VGND VGND VPWR VPWR _03597_ sky130_fd_sc_hd__o21ai_2
X_13004_ _04975_ _05508_ VGND VGND VPWR VPWR _05509_ sky130_fd_sc_hd__or2_2
X_10216_ _02125_ _02128_ _02124_ VGND VGND VPWR VPWR _02446_ sky130_fd_sc_hd__a21o_1
XFILLER_0_120_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11196_ _03520_ _03240_ VGND VGND VPWR VPWR _03522_ sky130_fd_sc_hd__nor2_1
XANTENNA__11547__D _02120_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10147_ _02366_ _04048_ _05027_ _02369_ VGND VGND VPWR VPWR _02370_ sky130_fd_sc_hd__and4b_1
XFILLER_0_118_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10078_ _02282_ _02293_ VGND VGND VPWR VPWR _02294_ sky130_fd_sc_hd__and2_1
X_13906_ _06413_ _06386_ _06411_ VGND VGND VPWR VPWR _06484_ sky130_fd_sc_hd__nor3_1
XANTENNA__07688__A2 _03499_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12681__A2 _05150_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07115__A _00563_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13837_ _06405_ _06407_ VGND VGND VPWR VPWR _06408_ sky130_fd_sc_hd__nand2_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10179__C _06744_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13768_ _05867_ _05882_ VGND VGND VPWR VPWR _06332_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12719_ _05193_ _05195_ VGND VGND VPWR VPWR _05196_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_17_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10476__A _02728_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13699_ _06254_ _06255_ _02427_ _02720_ VGND VGND VPWR VPWR _06256_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_26_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09930_ _02130_ _02131_ VGND VGND VPWR VPWR _02132_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09861_ _02031_ _02033_ VGND VGND VPWR VPWR _02056_ sky130_fd_sc_hd__nor2_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08812_ _00906_ _00907_ VGND VGND VPWR VPWR _00908_ sky130_fd_sc_hd__xor2_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09792_ _01792_ _01793_ VGND VGND VPWR VPWR _01981_ sky130_fd_sc_hd__nor2_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09505__A _02116_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08743_ _00824_ _00832_ VGND VGND VPWR VPWR _00833_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08674_ _00754_ _00756_ VGND VGND VPWR VPWR _00757_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07625_ _05467_ _00541_ VGND VGND VPWR VPWR _06208_ sky130_fd_sc_hd__nand2_1
XTAP_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12866__A _02008_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11770__A _05445_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07556_ _03147_ VGND VGND VPWR VPWR _05467_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_76_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07487_ _04697_ _04675_ VGND VGND VPWR VPWR _04708_ sky130_fd_sc_hd__and2b_1
XFILLER_0_63_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09226_ _00410_ _00376_ _00380_ _03015_ VGND VGND VPWR VPWR _01362_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_119_788 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13697__A _00416_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09157_ _01221_ _01283_ VGND VGND VPWR VPWR _01286_ sky130_fd_sc_hd__nand2_1
XANTENNA__09894__B _06450_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10738__A2 _02758_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08108_ _05478_ _00094_ VGND VGND VPWR VPWR _00152_ sky130_fd_sc_hd__nand2_1
X_09088_ net16 VGND VGND VPWR VPWR _01211_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_31_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08039_ _00081_ _07077_ _00082_ VGND VGND VPWR VPWR _00083_ sky130_fd_sc_hd__and3_1
XFILLER_0_101_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11050_ _03355_ _03358_ _03360_ VGND VGND VPWR VPWR _03361_ sky130_fd_sc_hd__o21a_1
XANTENNA__08564__B1 _00526_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10001_ _01869_ _01885_ _01887_ VGND VGND VPWR VPWR _02210_ sky130_fd_sc_hd__a21bo_1
XANTENNA__13582__D _03783_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11952_ _04349_ _04350_ VGND VGND VPWR VPWR _04352_ sky130_fd_sc_hd__and2_1
X_10903_ _03197_ _03198_ VGND VGND VPWR VPWR _03199_ sky130_fd_sc_hd__nor2_1
X_11883_ _04072_ _04096_ _04098_ _04275_ VGND VGND VPWR VPWR _04276_ sky130_fd_sc_hd__a211o_1
XFILLER_0_98_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13622_ _06017_ _06030_ VGND VGND VPWR VPWR _06171_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10834_ _03111_ _03115_ VGND VGND VPWR VPWR _03123_ sky130_fd_sc_hd__xor2_1
XFILLER_0_13_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12495__B _03938_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13553_ _06092_ _06068_ _06094_ VGND VGND VPWR VPWR _06095_ sky130_fd_sc_hd__nor3_1
XFILLER_0_137_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__07589__B _05467_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10765_ _01156_ _02766_ _02998_ _02999_ VGND VGND VPWR VPWR _03047_ sky130_fd_sc_hd__a211o_1
XFILLER_0_66_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12504_ _04946_ _04945_ VGND VGND VPWR VPWR _04959_ sky130_fd_sc_hd__or2b_1
XFILLER_0_81_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13484_ _06009_ _06018_ _01957_ _03690_ VGND VGND VPWR VPWR _06019_ sky130_fd_sc_hd__and4_1
X_10696_ _02955_ _02952_ VGND VGND VPWR VPWR _02972_ sky130_fd_sc_hd__xor2_1
XFILLER_0_125_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12435_ _04826_ _04882_ VGND VGND VPWR VPWR _04883_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_745 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12366_ _04805_ _04804_ VGND VGND VPWR VPWR _04808_ sky130_fd_sc_hd__or2b_1
XFILLER_0_23_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14105_ _06666_ _06670_ _06668_ VGND VGND VPWR VPWR _06700_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_1_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11317_ _02796_ _02918_ VGND VGND VPWR VPWR _03655_ sky130_fd_sc_hd__nor2_1
XFILLER_0_50_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09309__B _00818_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12297_ _04729_ _04731_ VGND VGND VPWR VPWR _04732_ sky130_fd_sc_hd__nor2_1
X_14036_ _06492_ _06625_ VGND VGND VPWR VPWR _06627_ sky130_fd_sc_hd__xor2_4
XANTENNA_output75_A net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09347__A2 _04015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11248_ _03562_ _03563_ VGND VGND VPWR VPWR _03579_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07358__A1 _01295_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07358__B2 _01306_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12351__B2 _03696_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11179_ _03402_ _03441_ _03386_ VGND VGND VPWR VPWR _03503_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_38_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07771__C _04851_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_244 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12654__A2 _02759_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07410_ _03850_ _01394_ net8 _03718_ VGND VGND VPWR VPWR _03861_ sky130_fd_sc_hd__and4_1
XFILLER_0_9_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08390_ _00445_ _00446_ VGND VGND VPWR VPWR _00447_ sky130_fd_sc_hd__and2b_1
XANTENNA__12406__A2 _00413_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09060__A _01179_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07341_ _03092_ VGND VGND VPWR VPWR _03103_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07272_ _00453_ _02335_ _02313_ VGND VGND VPWR VPWR _02346_ sky130_fd_sc_hd__a21o_1
XFILLER_0_116_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09011_ _00003_ _00151_ VGND VGND VPWR VPWR _01126_ sky130_fd_sc_hd__nand2_1
XFILLER_0_143_544 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11393__A2 _01179_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09913_ _02007_ _02040_ _01179_ _01254_ VGND VGND VPWR VPWR _02113_ sky130_fd_sc_hd__nand4_2
XANTENNA__12342__A1 _01260_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11765__A _02280_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07962__B _02171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09844_ _01825_ _01827_ _02034_ VGND VGND VPWR VPWR _02038_ sky130_fd_sc_hd__and3_2
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09235__A _01284_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07681__C net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09775_ _01813_ _01816_ VGND VGND VPWR VPWR _01962_ sky130_fd_sc_hd__and2_1
X_08726_ _00640_ _00812_ VGND VGND VPWR VPWR _00815_ sky130_fd_sc_hd__nand2_1
XTAP_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08657_ _00578_ _00736_ VGND VGND VPWR VPWR _00739_ sky130_fd_sc_hd__nand2_1
XANTENNA__12596__A _00745_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07608_ _03103_ _05800_ VGND VGND VPWR VPWR _06021_ sky130_fd_sc_hd__nand2_1
XTAP_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08588_ _00634_ _00663_ VGND VGND VPWR VPWR _00664_ sky130_fd_sc_hd__nor2_1
XANTENNA__11931__C _00572_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10828__B _02724_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07539_ _05170_ _05269_ VGND VGND VPWR VPWR _05280_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10959__A2 _01400_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10547__C _02725_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07202__B _00300_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10550_ _02808_ _02809_ _02807_ VGND VGND VPWR VPWR _02811_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_107_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07824__A2 net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09209_ _01341_ _01342_ VGND VGND VPWR VPWR _01343_ sky130_fd_sc_hd__nor2_1
X_10481_ _02726_ VGND VGND VPWR VPWR _02735_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_106_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12220_ _04645_ _04646_ VGND VGND VPWR VPWR _04647_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13577__D _02857_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12581__A1 _00742_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12151_ _04568_ _04563_ _04569_ VGND VGND VPWR VPWR _04571_ sky130_fd_sc_hd__nand3_2
XANTENNA__12581__B2 _00392_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09129__B _00322_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11102_ _03412_ _03417_ VGND VGND VPWR VPWR _03418_ sky130_fd_sc_hd__nor2_2
X_12082_ _04413_ _04493_ VGND VGND VPWR VPWR _04495_ sky130_fd_sc_hd__nor2_1
X_11033_ _03338_ _03341_ VGND VGND VPWR VPWR _03342_ sky130_fd_sc_hd__nor2_1
XANTENNA__07872__B _00410_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09145__A net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07760__A1 _00442_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12984_ _05450_ _05486_ VGND VGND VPWR VPWR _05487_ sky130_fd_sc_hd__nor2_2
XFILLER_0_99_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11935_ _00003_ _01585_ _04332_ VGND VGND VPWR VPWR _04333_ sky130_fd_sc_hd__and3_1
XANTENNA_output113_A net129 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11866_ _00113_ _00258_ _00415_ _00574_ VGND VGND VPWR VPWR _04258_ sky130_fd_sc_hd__and4_1
XFILLER_0_86_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13597__B1 _02856_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13605_ _06147_ net141 _06151_ VGND VGND VPWR VPWR _06152_ sky130_fd_sc_hd__o21a_1
XFILLER_0_145_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10817_ _03068_ _03104_ VGND VGND VPWR VPWR _03105_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_138_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_848 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11797_ _04173_ _04175_ _04179_ _04181_ VGND VGND VPWR VPWR _04182_ sky130_fd_sc_hd__o211a_1
XFILLER_0_131_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13536_ _02722_ VGND VGND VPWR VPWR _06077_ sky130_fd_sc_hd__buf_2
XFILLER_0_55_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10748_ _03025_ _03028_ VGND VGND VPWR VPWR _03029_ sky130_fd_sc_hd__and2_1
XFILLER_0_137_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13467_ _05998_ _06000_ VGND VGND VPWR VPWR _06001_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_70_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10679_ _02982_ _01546_ _02156_ _00377_ VGND VGND VPWR VPWR _02953_ sky130_fd_sc_hd__a22o_1
XANTENNA__10754__A _00399_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12418_ _00375_ _00378_ _00414_ _00572_ VGND VGND VPWR VPWR _04865_ sky130_fd_sc_hd__and4_2
XFILLER_0_106_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13398_ _05914_ _05395_ _05924_ VGND VGND VPWR VPWR _05926_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08224__A _00101_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10032__C1 _01867_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12349_ _01260_ _00605_ VGND VGND VPWR VPWR _04789_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14019_ _06491_ _06504_ VGND VGND VPWR VPWR _06608_ sky130_fd_sc_hd__nor2_1
X_07890_ _02719_ _00475_ _06945_ VGND VGND VPWR VPWR _07019_ sky130_fd_sc_hd__and3_1
XFILLER_0_65_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09560_ _00654_ _01472_ _01724_ _01725_ VGND VGND VPWR VPWR _01727_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_65_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08511_ _00576_ _00578_ VGND VGND VPWR VPWR _00579_ sky130_fd_sc_hd__and2_1
X_09491_ _00431_ _04169_ net51 net52 VGND VGND VPWR VPWR _01651_ sky130_fd_sc_hd__and4_1
XFILLER_0_77_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08442_ _00502_ _00503_ VGND VGND VPWR VPWR _00504_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_247 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08373_ _00421_ _00427_ VGND VGND VPWR VPWR _00428_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_135_308 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07324_ _02894_ _02905_ VGND VGND VPWR VPWR _02916_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07255_ _02149_ VGND VGND VPWR VPWR _02160_ sky130_fd_sc_hd__buf_2
XANTENNA__09008__A1 _03004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09008__B2 _00095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13040__A _05536_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_143_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07186_ _01394_ VGND VGND VPWR VPWR _01405_ sky130_fd_sc_hd__buf_4
XANTENNA__08134__A _00100_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13512__B1 _02737_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09827_ _02012_ _02019_ VGND VGND VPWR VPWR _02020_ sky130_fd_sc_hd__xor2_1
X_09758_ _01663_ _01696_ _01943_ VGND VGND VPWR VPWR _01944_ sky130_fd_sc_hd__a21o_1
XANTENNA__07526__A1_N _00901_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08709_ _00794_ _00795_ VGND VGND VPWR VPWR _00796_ sky130_fd_sc_hd__xnor2_1
XTAP_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09689_ _01754_ _01867_ VGND VGND VPWR VPWR _01868_ sky130_fd_sc_hd__xnor2_2
XTAP_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11720_ _04072_ _04096_ VGND VGND VPWR VPWR _04097_ sky130_fd_sc_hd__xor2_1
XFILLER_0_96_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10558__B _02169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11651_ _03844_ _04012_ _04020_ VGND VGND VPWR VPWR _04021_ sky130_fd_sc_hd__a21oi_1
XTAP_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10602_ _02866_ _02867_ _00142_ _01059_ VGND VGND VPWR VPWR _02868_ sky130_fd_sc_hd__and4b_1
XFILLER_0_36_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11582_ _03830_ _03831_ VGND VGND VPWR VPWR _03945_ sky130_fd_sc_hd__or2_1
XFILLER_0_52_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13321_ _05647_ _05663_ _05826_ VGND VGND VPWR VPWR _05842_ sky130_fd_sc_hd__nand3_2
XFILLER_0_107_544 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10533_ _02746_ _02790_ _02791_ VGND VGND VPWR VPWR _02792_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_134_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12492__C _03685_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13252_ _05546_ _05777_ VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__xnor2_2
XFILLER_0_107_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10464_ _02274_ _02276_ _02491_ _02715_ _02716_ VGND VGND VPWR VPWR _02717_ sky130_fd_sc_hd__a32o_1
XFILLER_0_51_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12203_ _04626_ _04627_ VGND VGND VPWR VPWR _04628_ sky130_fd_sc_hd__or2_1
XFILLER_0_32_372 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13183_ _05685_ _05688_ VGND VGND VPWR VPWR _05706_ sky130_fd_sc_hd__xor2_4
X_10395_ _02392_ _02421_ VGND VGND VPWR VPWR _02641_ sky130_fd_sc_hd__and2_1
XANTENNA__08979__A _03268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12134_ _04546_ _04551_ VGND VGND VPWR VPWR _04552_ sky130_fd_sc_hd__or2b_1
XANTENNA__07883__A net177 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09970__A2 _01060_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12065_ _04247_ _04249_ VGND VGND VPWR VPWR _04476_ sky130_fd_sc_hd__xor2_1
XFILLER_0_19_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11016_ _02552_ _02556_ _03322_ VGND VGND VPWR VPWR _03324_ sky130_fd_sc_hd__a21o_1
XFILLER_0_126_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12948__B _05447_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__14074__A4 _02743_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12967_ _05468_ VGND VGND VPWR VPWR _05469_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11918_ _04313_ _04314_ VGND VGND VPWR VPWR _04315_ sky130_fd_sc_hd__or2b_1
XANTENNA__10096__A2 net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12898_ _05383_ _05392_ VGND VGND VPWR VPWR _05393_ sky130_fd_sc_hd__xor2_1
XANTENNA__08219__A _06966_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07123__A net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12386__D _00734_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11849_ _04219_ _04222_ VGND VGND VPWR VPWR _04239_ sky130_fd_sc_hd__and2_1
XFILLER_0_74_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10187__C net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09789__A2 _01181_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12793__A1 _02728_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13519_ _06055_ _06056_ VGND VGND VPWR VPWR _06058_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_188 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07777__B net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10484__A _01473_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11348__A2 _01956_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13010__D _05515_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08889__A _06965_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08991_ _01102_ _01103_ VGND VGND VPWR VPWR _01104_ sky130_fd_sc_hd__and2b_1
X_07942_ _07069_ _07070_ VGND VGND VPWR VPWR _07071_ sky130_fd_sc_hd__nor2_1
X_07873_ _06975_ _06973_ VGND VGND VPWR VPWR _07002_ sky130_fd_sc_hd__and2b_1
XANTENNA__07724__A1 _02259_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07724__B2 _02171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09612_ _01779_ _01782_ _01783_ VGND VGND VPWR VPWR _01784_ sky130_fd_sc_hd__nor3_1
XFILLER_0_92_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09543_ _01703_ _01707_ VGND VGND VPWR VPWR _01708_ sky130_fd_sc_hd__xor2_1
XANTENNA__11762__B _02018_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12577__C _01934_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09474_ _01439_ _01631_ _01632_ _01428_ VGND VGND VPWR VPWR _01633_ sky130_fd_sc_hd__or4b_4
X_08425_ _00260_ _00265_ _00483_ VGND VGND VPWR VPWR _00485_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_46_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11036__A1 _00142_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08356_ _00400_ _00406_ _00408_ _00409_ VGND VGND VPWR VPWR _00411_ sky130_fd_sc_hd__a31o_2
XANTENNA__11036__B2 _00778_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07307_ _01470_ _02719_ VGND VGND VPWR VPWR _02729_ sky130_fd_sc_hd__nand2_1
X_08287_ _00332_ _00334_ VGND VGND VPWR VPWR _00335_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_116_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07238_ _01930_ _01963_ VGND VGND VPWR VPWR _01974_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07169_ _00880_ net26 _01197_ _01208_ VGND VGND VPWR VPWR _01219_ sky130_fd_sc_hd__and4_1
XFILLER_0_30_854 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_720 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10180_ _02404_ _02405_ VGND VGND VPWR VPWR _02406_ sky130_fd_sc_hd__or2_1
XFILLER_0_100_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07208__A _00891_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13870_ _06431_ _06443_ VGND VGND VPWR VPWR _06444_ sky130_fd_sc_hd__or2_1
X_12821_ _05039_ _05130_ VGND VGND VPWR VPWR _05308_ sky130_fd_sc_hd__nand2_1
XANTENNA__13590__D _02858_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12752_ _05230_ _05231_ VGND VGND VPWR VPWR _05232_ sky130_fd_sc_hd__or2_1
XTAP_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10288__B _05742_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11703_ _04076_ _02627_ _04077_ VGND VGND VPWR VPWR _04078_ sky130_fd_sc_hd__and3_1
XTAP_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12683_ _05141_ _05142_ _05144_ VGND VGND VPWR VPWR _05156_ sky130_fd_sc_hd__o21a_1
XTAP_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12784__A _00414_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11027__A1 _05027_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11634_ _03956_ _04001_ VGND VGND VPWR VPWR _04002_ sky130_fd_sc_hd__nor2_1
XANTENNA__07878__A _01230_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11027__B2 _04851_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11565_ _00486_ _02117_ VGND VGND VPWR VPWR _03926_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13304_ _05678_ _05825_ VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__xor2_2
XFILLER_0_122_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10516_ _02771_ _02772_ VGND VGND VPWR VPWR _02774_ sky130_fd_sc_hd__or2b_1
XFILLER_0_134_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11496_ _03789_ _03838_ _03790_ _03800_ VGND VGND VPWR VPWR _03851_ sky130_fd_sc_hd__or4_1
XFILLER_0_12_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_810 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13235_ _05575_ _05579_ _05585_ _05591_ _05589_ VGND VGND VPWR VPWR _05760_ sky130_fd_sc_hd__a32o_1
X_10447_ _02694_ _02698_ VGND VGND VPWR VPWR _02699_ sky130_fd_sc_hd__xnor2_2
XANTENNA__10538__B1 _02728_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13166_ _04546_ _05686_ VGND VGND VPWR VPWR _05688_ sky130_fd_sc_hd__xnor2_4
X_10378_ _02621_ _02622_ VGND VGND VPWR VPWR _02623_ sky130_fd_sc_hd__xor2_1
X_12117_ _04492_ _04533_ VGND VGND VPWR VPWR _04534_ sky130_fd_sc_hd__xnor2_4
X_13097_ _04592_ _04588_ _05611_ VGND VGND VPWR VPWR _05612_ sky130_fd_sc_hd__o21a_1
XANTENNA__07118__A net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12048_ _04142_ _04252_ VGND VGND VPWR VPWR _04458_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_137_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10479__A _01472_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13999_ _06562_ _06585_ VGND VGND VPWR VPWR _06586_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_854 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08210_ _00137_ _00175_ VGND VGND VPWR VPWR _00254_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09190_ _01320_ _01321_ VGND VGND VPWR VPWR _01322_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10926__B _02758_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08141_ _06985_ _07082_ VGND VGND VPWR VPWR _00185_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08072_ _01350_ _00113_ _00115_ VGND VGND VPWR VPWR _00116_ sky130_fd_sc_hd__and3_1
XFILLER_0_113_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09934__A2 _01954_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08974_ _00949_ _00952_ _01084_ VGND VGND VPWR VPWR _01085_ sky130_fd_sc_hd__o21a_1
XANTENNA__09227__B _02960_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11476__C _01954_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07925_ _07052_ _07053_ VGND VGND VPWR VPWR _07054_ sky130_fd_sc_hd__and2b_1
X_07856_ _06899_ _06984_ VGND VGND VPWR VPWR _06985_ sky130_fd_sc_hd__and2b_1
XANTENNA__07173__A2 _00672_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07787_ _06914_ _06915_ VGND VGND VPWR VPWR _06916_ sky130_fd_sc_hd__xnor2_1
X_09526_ _01686_ _01688_ VGND VGND VPWR VPWR _01690_ sky130_fd_sc_hd__and2b_1
XFILLER_0_79_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09457_ _06820_ net8 net9 net64 VGND VGND VPWR VPWR _01615_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08408_ _00283_ _00284_ VGND VGND VPWR VPWR _00467_ sky130_fd_sc_hd__nand2_1
XANTENNA__11009__A1 _05203_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11009__B2 _01369_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12206__B1 _02134_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09388_ _01529_ _01538_ VGND VGND VPWR VPWR _01539_ sky130_fd_sc_hd__xnor2_2
XANTENNA__10480__A2 _02722_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10836__B _01933_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08339_ _03740_ VGND VGND VPWR VPWR _00392_ sky130_fd_sc_hd__buf_4
XANTENNA__10555__C _00095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11350_ _03687_ VGND VGND VPWR VPWR _03690_ sky130_fd_sc_hd__buf_2
XFILLER_0_117_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10301_ _02504_ _02537_ VGND VGND VPWR VPWR _02538_ sky130_fd_sc_hd__xnor2_2
XANTENNA__13706__B1 _02725_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11281_ _03613_ _03614_ VGND VGND VPWR VPWR _03615_ sky130_fd_sc_hd__nand2_1
XFILLER_0_132_686 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13020_ _01637_ net131 _01433_ _02046_ VGND VGND VPWR VPWR _05527_ sky130_fd_sc_hd__and4_1
X_10232_ _00322_ _02459_ _02461_ _02462_ VGND VGND VPWR VPWR _02463_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__11667__B _06885_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08322__A _04015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10571__B _03015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10163_ _02385_ _02386_ VGND VGND VPWR VPWR _02387_ sky130_fd_sc_hd__nand2_1
X_10094_ _02309_ _02310_ VGND VGND VPWR VPWR _02311_ sky130_fd_sc_hd__xnor2_2
XANTENNA__13485__A2 _01957_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08976__B net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13922_ _06499_ _06500_ VGND VGND VPWR VPWR _06501_ sky130_fd_sc_hd__and2_1
XFILLER_0_16_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13853_ _01517_ _03679_ _05386_ VGND VGND VPWR VPWR _06425_ sky130_fd_sc_hd__and3_1
XFILLER_0_69_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12804_ _05056_ _05110_ VGND VGND VPWR VPWR _05289_ sky130_fd_sc_hd__nand2_1
X_10996_ _03265_ _03300_ VGND VGND VPWR VPWR _03302_ sky130_fd_sc_hd__xnor2_1
X_13784_ _05891_ _05894_ VGND VGND VPWR VPWR _06349_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12735_ _05145_ _05150_ _05153_ VGND VGND VPWR VPWR _05213_ sky130_fd_sc_hd__o21ai_1
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08664__A2 _00745_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12666_ _05133_ _05134_ _05136_ VGND VGND VPWR VPWR _05138_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_72_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14218__B _00344_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07401__A net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11617_ _03981_ _03973_ VGND VGND VPWR VPWR _03984_ sky130_fd_sc_hd__xor2_4
XFILLER_0_65_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12597_ _03740_ _01411_ _02849_ _03707_ VGND VGND VPWR VPWR _05062_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07120__B _00650_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11548_ _06964_ _02119_ _02120_ _00121_ VGND VGND VPWR VPWR _03908_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11479_ _03830_ _03831_ VGND VGND VPWR VPWR _03832_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13218_ _05667_ _05677_ VGND VGND VPWR VPWR _05745_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09328__A _01472_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14198_ _06622_ _06791_ VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__xor2_4
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13149_ _03053_ _04624_ VGND VGND VPWR VPWR _05669_ sky130_fd_sc_hd__xnor2_2
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11296__C _02736_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07710_ _06836_ _06838_ VGND VGND VPWR VPWR _06839_ sky130_fd_sc_hd__and2b_1
X_08690_ _00773_ _00774_ VGND VGND VPWR VPWR _00775_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09063__A _01182_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07641_ _06362_ _06373_ VGND VGND VPWR VPWR _06384_ sky130_fd_sc_hd__nor2_1
XANTENNA__12839__D _02727_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07572_ _05555_ _05610_ _03301_ VGND VGND VPWR VPWR _05643_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_76_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09311_ _01449_ _01327_ _01453_ VGND VGND VPWR VPWR _01454_ sky130_fd_sc_hd__nor3_1
XFILLER_0_48_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09242_ _01366_ _01081_ _01377_ VGND VGND VPWR VPWR _01379_ sky130_fd_sc_hd__nor3_1
XFILLER_0_29_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09510__B _00458_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_255 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09173_ _01301_ _01302_ VGND VGND VPWR VPWR _01303_ sky130_fd_sc_hd__nand2_1
XANTENNA__12209__A2_N _03682_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08124_ _00166_ _00167_ VGND VGND VPWR VPWR _00168_ sky130_fd_sc_hd__nor2_1
XANTENNA__11962__A2 _03678_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08055_ _00000_ _00097_ VGND VGND VPWR VPWR _00099_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13686__C _02735_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12590__C _02855_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10822__D net57 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08957_ _02467_ _01066_ VGND VGND VPWR VPWR _01067_ sky130_fd_sc_hd__nand2_1
X_07908_ _07003_ _07036_ VGND VGND VPWR VPWR _07037_ sky130_fd_sc_hd__xor2_1
X_08888_ _00806_ _00837_ VGND VGND VPWR VPWR _00992_ sky130_fd_sc_hd__or2b_1
XANTENNA__12675__B1 _00381_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07839_ _06824_ _06877_ VGND VGND VPWR VPWR _06968_ sky130_fd_sc_hd__and2_1
XANTENNA__11008__A _00294_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10850_ _05566_ _01410_ _03139_ _03140_ VGND VGND VPWR VPWR _03141_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_67_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09509_ _01532_ _01533_ _01531_ VGND VGND VPWR VPWR _01671_ sky130_fd_sc_hd__o21ai_1
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_846 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10781_ _06937_ _06494_ _02725_ _02730_ VGND VGND VPWR VPWR _03065_ sky130_fd_sc_hd__and4_1
XFILLER_0_39_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12520_ _04967_ _04975_ _04976_ VGND VGND VPWR VPWR _04977_ sky130_fd_sc_hd__a21oi_2
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12451_ _04871_ _04847_ VGND VGND VPWR VPWR _04901_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11402_ _03736_ _03739_ _03746_ VGND VGND VPWR VPWR _03747_ sky130_fd_sc_hd__o21ai_2
X_12382_ _04783_ _04786_ VGND VGND VPWR VPWR _04825_ sky130_fd_sc_hd__xor2_1
XFILLER_0_117_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14121_ _06657_ _06717_ VGND VGND VPWR VPWR _06718_ sky130_fd_sc_hd__nand2_1
X_11333_ _03669_ _03671_ VGND VGND VPWR VPWR _03672_ sky130_fd_sc_hd__nand2_1
XFILLER_0_132_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10582__A _00310_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14052_ _06635_ _06643_ VGND VGND VPWR VPWR _06644_ sky130_fd_sc_hd__or2_1
X_11264_ _03591_ _03592_ VGND VGND VPWR VPWR _03596_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08052__A _00497_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13003_ _04973_ _04974_ VGND VGND VPWR VPWR _05508_ sky130_fd_sc_hd__nor2_1
X_10215_ _02442_ _02443_ VGND VGND VPWR VPWR _02444_ sky130_fd_sc_hd__nor2_1
X_11195_ _03192_ _03199_ _03204_ VGND VGND VPWR VPWR _03520_ sky130_fd_sc_hd__nor3_1
X_10146_ _04851_ _04015_ _00780_ net4 VGND VGND VPWR VPWR _02369_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10077_ _02290_ _02292_ VGND VGND VPWR VPWR _02293_ sky130_fd_sc_hd__and2b_1
XFILLER_0_27_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12302__A _00415_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13905_ _06451_ _06479_ _06481_ VGND VGND VPWR VPWR _06482_ sky130_fd_sc_hd__o21a_1
XFILLER_0_134_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13836_ _06397_ _06402_ _06404_ VGND VGND VPWR VPWR _06407_ sky130_fd_sc_hd__or3_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12956__B _05429_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10979_ _03271_ _03274_ VGND VGND VPWR VPWR _03283_ sky130_fd_sc_hd__or2_1
X_13767_ _06328_ _06330_ VGND VGND VPWR VPWR _06331_ sky130_fd_sc_hd__nor2_1
XANTENNA__14229__A _06810_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12718_ _05178_ _05194_ VGND VGND VPWR VPWR _05195_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_84_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13698_ _01289_ _02726_ _02730_ _01188_ VGND VGND VPWR VPWR _06255_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_38_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12972__A _05451_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12649_ _02008_ _01061_ VGND VGND VPWR VPWR _05119_ sky130_fd_sc_hd__nand2_1
XFILLER_0_111_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_472 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09058__A _01177_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09860_ _02053_ _02039_ _02054_ VGND VGND VPWR VPWR _02055_ sky130_fd_sc_hd__a21o_2
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08811_ _00300_ net16 VGND VGND VPWR VPWR _00907_ sky130_fd_sc_hd__and2_1
X_09791_ _01959_ _01979_ VGND VGND VPWR VPWR _01980_ sky130_fd_sc_hd__xnor2_2
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08742_ _00830_ _00831_ VGND VGND VPWR VPWR _00832_ sky130_fd_sc_hd__or2_1
XANTENNA__07306__A net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08673_ _02029_ _00755_ VGND VGND VPWR VPWR _00756_ sky130_fd_sc_hd__nand2_1
XFILLER_0_108_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07624_ _05445_ _05467_ _05742_ _02664_ VGND VGND VPWR VPWR _06197_ sky130_fd_sc_hd__and4_1
XTAP_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12866__B _02765_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07555_ _05445_ VGND VGND VPWR VPWR _05456_ sky130_fd_sc_hd__buf_4
XANTENNA__11770__B _05731_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07486_ _04631_ _04686_ VGND VGND VPWR VPWR _04697_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09225_ _01057_ _01107_ _01110_ VGND VGND VPWR VPWR _01360_ sky130_fd_sc_hd__o21a_1
XFILLER_0_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09156_ _01221_ _01283_ VGND VGND VPWR VPWR _01285_ sky130_fd_sc_hd__or2_1
XANTENNA__13697__B _01288_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09894__C _02090_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08107_ _05181_ VGND VGND VPWR VPWR _00151_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_32_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09087_ _03850_ _00730_ net15 _01306_ VGND VGND VPWR VPWR _01210_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_142_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08038_ _00041_ _00042_ _00078_ _00079_ VGND VGND VPWR VPWR _00082_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_101_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10000_ _02184_ _02208_ VGND VGND VPWR VPWR _02209_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08564__A1 _00519_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08564__B2 _03554_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09989_ _02195_ _02196_ VGND VGND VPWR VPWR _02197_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11951_ _04349_ _04350_ VGND VGND VPWR VPWR _04351_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11961__A _03059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10902_ _03178_ _03181_ VGND VGND VPWR VPWR _03198_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11882_ _00262_ _00263_ _02090_ _01780_ VGND VGND VPWR VPWR _04275_ sky130_fd_sc_hd__and4_1
XFILLER_0_67_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09431__A _01272_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13621_ _06119_ _06130_ _06168_ _06118_ VGND VGND VPWR VPWR _06170_ sky130_fd_sc_hd__o31ai_1
X_10833_ _03120_ _03121_ VGND VGND VPWR VPWR _03122_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_67_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13552_ _06062_ _06093_ VGND VGND VPWR VPWR _06094_ sky130_fd_sc_hd__xor2_1
XFILLER_0_67_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10764_ _02998_ _02999_ _01156_ _02766_ VGND VGND VPWR VPWR _03046_ sky130_fd_sc_hd__o211ai_1
XANTENNA__07589__C _02105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08047__A _03521_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12503_ _00378_ _00741_ _04957_ VGND VGND VPWR VPWR _04958_ sky130_fd_sc_hd__and3_1
X_13483_ _02858_ VGND VGND VPWR VPWR _06018_ sky130_fd_sc_hd__buf_2
XFILLER_0_54_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10695_ _02968_ _02969_ VGND VGND VPWR VPWR _02970_ sky130_fd_sc_hd__nand2_1
XFILLER_0_109_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13376__A1 _00607_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12434_ _04825_ _04798_ _04824_ VGND VGND VPWR VPWR _04882_ sky130_fd_sc_hd__or3_1
XFILLER_0_35_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12365_ _04804_ _04805_ VGND VGND VPWR VPWR _04806_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_105_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14104_ _06644_ _06697_ _06698_ VGND VGND VPWR VPWR _06699_ sky130_fd_sc_hd__or3_4
X_11316_ _03651_ _03652_ VGND VGND VPWR VPWR _03654_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12296_ _02427_ _02190_ _02088_ _02188_ VGND VGND VPWR VPWR _04731_ sky130_fd_sc_hd__a22oi_1
X_14035_ _06624_ _06607_ _06506_ VGND VGND VPWR VPWR _06625_ sky130_fd_sc_hd__a21o_1
XFILLER_0_129_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11247_ _03575_ _03577_ VGND VGND VPWR VPWR _03578_ sky130_fd_sc_hd__or2_1
XANTENNA__07358__A2 _02664_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09606__A _03059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11178_ _03205_ _03242_ _03189_ VGND VGND VPWR VPWR _03502_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10362__A1 _06744_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10129_ _02212_ _02216_ VGND VGND VPWR VPWR _02350_ sky130_fd_sc_hd__and2_1
XANTENNA__07771__D net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09504__B1 _01505_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13819_ _02187_ _01955_ _03686_ _01400_ VGND VGND VPWR VPWR _06388_ sky130_fd_sc_hd__a22o_1
XANTENNA__10487__A _02737_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07340_ _02007_ _02029_ _02105_ _02149_ VGND VGND VPWR VPWR _03092_ sky130_fd_sc_hd__and4_1
XFILLER_0_85_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_484 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07271_ _02280_ VGND VGND VPWR VPWR _02335_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__13798__A _02188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09010_ _01123_ _01124_ VGND VGND VPWR VPWR _01125_ sky130_fd_sc_hd__nor2_1
XFILLER_0_115_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_543 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09912_ _03070_ _01180_ _01249_ _02335_ VGND VGND VPWR VPWR _02112_ sky130_fd_sc_hd__a22o_1
XANTENNA__10950__A _00143_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12342__A2 _00605_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09843_ _02035_ _02034_ VGND VGND VPWR VPWR _02037_ sky130_fd_sc_hd__and2_2
XANTENNA__11765__B _03682_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07962__C _00004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09235__B _01230_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09774_ _00322_ _01960_ _01814_ VGND VGND VPWR VPWR _01961_ sky130_fd_sc_hd__and3_1
XANTENNA__07681__D net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08725_ _00640_ _00812_ VGND VGND VPWR VPWR _00813_ sky130_fd_sc_hd__or2_1
XTAP_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12877__A _01507_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08656_ _00578_ _00736_ VGND VGND VPWR VPWR _00738_ sky130_fd_sc_hd__or2_1
XTAP_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12596__B _01059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07607_ _05676_ _05687_ VGND VGND VPWR VPWR _06010_ sky130_fd_sc_hd__xnor2_2
XTAP_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08587_ _00641_ _00662_ VGND VGND VPWR VPWR _00663_ sky130_fd_sc_hd__xnor2_1
XTAP_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11931__D _01272_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_440 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07538_ _05236_ _05258_ VGND VGND VPWR VPWR _05269_ sky130_fd_sc_hd__xor2_2
XFILLER_0_64_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10547__D _02730_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07469_ _00573_ VGND VGND VPWR VPWR _04510_ sky130_fd_sc_hd__buf_2
XFILLER_0_107_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09208_ _01144_ _01330_ _01340_ VGND VGND VPWR VPWR _01342_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10480_ _02247_ _02722_ _02732_ _02733_ VGND VGND VPWR VPWR _02734_ sky130_fd_sc_hd__a31o_1
XFILLER_0_91_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09139_ _01258_ _01265_ VGND VGND VPWR VPWR _01266_ sky130_fd_sc_hd__xor2_1
X_12150_ _04568_ _04569_ _04563_ VGND VGND VPWR VPWR _04570_ sky130_fd_sc_hd__a21o_1
XANTENNA__12581__A2 _02849_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09129__C _01179_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11101_ _03413_ _03416_ VGND VGND VPWR VPWR _03417_ sky130_fd_sc_hd__and2b_1
X_12081_ _04413_ _04493_ VGND VGND VPWR VPWR _04494_ sky130_fd_sc_hd__and2_1
X_11032_ _03339_ _03340_ VGND VGND VPWR VPWR _03341_ sky130_fd_sc_hd__or2_1
XANTENNA__11541__B1 _01564_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07760__A2 _06775_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12983_ _05024_ _05026_ VGND VGND VPWR VPWR _05486_ sky130_fd_sc_hd__and2_1
XFILLER_0_87_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11934_ _04329_ _04331_ VGND VGND VPWR VPWR _04332_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11865_ _04038_ _04039_ VGND VGND VPWR VPWR _04256_ sky130_fd_sc_hd__and2b_1
XANTENNA__13597__A1 _01413_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13604_ _06139_ _06135_ VGND VGND VPWR VPWR _06151_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10100__A _01933_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10816_ _06637_ _02731_ _03102_ VGND VGND VPWR VPWR _03104_ sky130_fd_sc_hd__and3_1
XANTENNA__13597__B2 _01180_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11796_ _01361_ _02459_ _02673_ _01405_ VGND VGND VPWR VPWR _04181_ sky130_fd_sc_hd__a22o_1
XFILLER_0_144_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13535_ _01958_ VGND VGND VPWR VPWR _06075_ sky130_fd_sc_hd__buf_2
XFILLER_0_131_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10747_ _03013_ _03027_ VGND VGND VPWR VPWR _03028_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_125_523 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13466_ _05985_ _02722_ VGND VGND VPWR VPWR _06000_ sky130_fd_sc_hd__nand2_1
X_10678_ _02950_ _02951_ VGND VGND VPWR VPWR _02952_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10754__B _02759_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08505__A _00571_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12417_ _04861_ _04863_ VGND VGND VPWR VPWR _04864_ sky130_fd_sc_hd__xnor2_4
X_13397_ _05914_ _05395_ _05924_ VGND VGND VPWR VPWR _05925_ sky130_fd_sc_hd__and3_1
XFILLER_0_112_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12348_ _04780_ _04779_ VGND VGND VPWR VPWR _04788_ sky130_fd_sc_hd__or2b_1
XFILLER_0_121_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11866__A _00113_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12279_ _04710_ _04701_ VGND VGND VPWR VPWR _04712_ sky130_fd_sc_hd__or2b_1
XFILLER_0_120_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14018_ _06598_ _06605_ _06606_ VGND VGND VPWR VPWR _06607_ sky130_fd_sc_hd__o21a_4
XFILLER_0_65_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08510_ _00577_ VGND VGND VPWR VPWR _00578_ sky130_fd_sc_hd__inv_2
X_09490_ _03587_ _01545_ net52 _03576_ VGND VGND VPWR VPWR _01650_ sky130_fd_sc_hd__a22oi_1
X_08441_ _03059_ _00158_ _00501_ VGND VGND VPWR VPWR _00503_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_147_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13588__A1 _01414_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11106__A _07040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07303__B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08372_ _00425_ _00426_ VGND VGND VPWR VPWR _00427_ sky130_fd_sc_hd__nor2_1
XFILLER_0_147_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_83 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07323_ _02445_ _02883_ VGND VGND VPWR VPWR _02905_ sky130_fd_sc_hd__or2_1
XFILLER_0_85_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07254_ _00650_ VGND VGND VPWR VPWR _02149_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_60_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09008__A2 _00113_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07185_ _01208_ VGND VGND VPWR VPWR _01394_ sky130_fd_sc_hd__buf_6
XFILLER_0_143_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11771__B1 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11776__A _05456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10680__A _00366_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10326__A1 _04851_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10326__B2 net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09826_ _02016_ _02017_ VGND VGND VPWR VPWR _02019_ sky130_fd_sc_hd__xnor2_1
X_09757_ _01663_ _01696_ _01712_ VGND VGND VPWR VPWR _01943_ sky130_fd_sc_hd__o21a_1
XTAP_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08708_ _04081_ net45 VGND VGND VPWR VPWR _00795_ sky130_fd_sc_hd__nand2_1
XTAP_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09688_ _01865_ _01866_ VGND VGND VPWR VPWR _01867_ sky130_fd_sc_hd__nor2_2
XFILLER_0_96_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08639_ _00718_ _00719_ VGND VGND VPWR VPWR _00720_ sky130_fd_sc_hd__xnor2_1
XTAP_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11650_ _04018_ _04019_ VGND VGND VPWR VPWR _04020_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10601_ _04862_ _01410_ _02158_ _04873_ VGND VGND VPWR VPWR _02867_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11581_ _03941_ _03942_ _03893_ VGND VGND VPWR VPWR _03944_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_64_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10855__A _06461_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10532_ _02741_ _02745_ _02738_ VGND VGND VPWR VPWR _02791_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_92_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13320_ _05647_ _05841_ VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__xor2_4
XFILLER_0_92_796 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12492__D _00423_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10463_ _02490_ VGND VGND VPWR VPWR _02716_ sky130_fd_sc_hd__inv_2
X_13251_ _05776_ _05773_ VGND VGND VPWR VPWR _05777_ sky130_fd_sc_hd__and2_4
XANTENNA__09076__A2_N net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_340 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12202_ _04024_ _04596_ VGND VGND VPWR VPWR _04627_ sky130_fd_sc_hd__xnor2_4
X_13182_ _05700_ _05704_ VGND VGND VPWR VPWR _05705_ sky130_fd_sc_hd__and2_2
X_10394_ _02638_ _02639_ VGND VGND VPWR VPWR _02640_ sky130_fd_sc_hd__or2_1
XFILLER_0_32_384 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12133_ _04548_ _04550_ VGND VGND VPWR VPWR _04551_ sky130_fd_sc_hd__xor2_4
XANTENNA__08979__B _04026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07883__B net149 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10590__A _02306_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12064_ _04137_ _04139_ VGND VGND VPWR VPWR _04475_ sky130_fd_sc_hd__xor2_1
X_11015_ _05181_ net45 _02553_ VGND VGND VPWR VPWR _03322_ sky130_fd_sc_hd__and3_1
XANTENNA__08995__A _01062_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12966_ _05464_ _05466_ VGND VGND VPWR VPWR _05468_ sky130_fd_sc_hd__xnor2_1
X_11917_ _04306_ _04311_ VGND VGND VPWR VPWR _04314_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12897_ _05384_ _05391_ VGND VGND VPWR VPWR _05392_ sky130_fd_sc_hd__xor2_1
XFILLER_0_142_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11848_ _02665_ _02682_ VGND VGND VPWR VPWR _04238_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10187__D _00730_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11779_ _04159_ _04160_ _04152_ _04154_ VGND VGND VPWR VPWR _04162_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_137_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10253__B1 _02151_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13518_ _06055_ _06056_ VGND VGND VPWR VPWR _06057_ sky130_fd_sc_hd__nor2_1
XANTENNA__10484__B _02247_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13449_ _05979_ _05980_ VGND VGND VPWR VPWR _05981_ sky130_fd_sc_hd__and2b_1
XFILLER_0_113_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08889__B _06966_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08990_ _01068_ _01101_ _01069_ VGND VGND VPWR VPWR _01103_ sky130_fd_sc_hd__or3_1
X_07941_ _07055_ _07068_ VGND VGND VPWR VPWR _07070_ sky130_fd_sc_hd__and2_1
X_07872_ _00530_ _00410_ VGND VGND VPWR VPWR _07001_ sky130_fd_sc_hd__nand2_1
XANTENNA__10005__A _05203_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07724__A2 _03543_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09611_ _02335_ _01780_ _01781_ VGND VGND VPWR VPWR _01783_ sky130_fd_sc_hd__a21oi_1
X_09542_ _01705_ _01706_ VGND VGND VPWR VPWR _01707_ sky130_fd_sc_hd__xor2_1
XFILLER_0_92_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11762__C _01953_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12577__D _02169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09473_ _01629_ _01630_ _01627_ _01628_ VGND VGND VPWR VPWR _01632_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_93_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08424_ _00483_ _00265_ _00260_ VGND VGND VPWR VPWR _00484_ sky130_fd_sc_hd__and3b_1
XFILLER_0_59_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_538 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08355_ _00387_ _00396_ _00398_ VGND VGND VPWR VPWR _00409_ sky130_fd_sc_hd__o21a_1
XANTENNA__11036__A2 _04037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07306_ net30 VGND VGND VPWR VPWR _02719_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_74_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08286_ _03532_ _00094_ VGND VGND VPWR VPWR _00334_ sky130_fd_sc_hd__nand2_1
XFILLER_0_117_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07237_ _01908_ _01919_ _01952_ VGND VGND VPWR VPWR _01963_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_15_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07168_ _00716_ VGND VGND VPWR VPWR _01208_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_131_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07099_ _00442_ VGND VGND VPWR VPWR _00453_ sky130_fd_sc_hd__buf_4
XFILLER_0_100_732 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07208__B _00672_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09704__A _00388_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09809_ _01791_ _01794_ _01999_ VGND VGND VPWR VPWR _02000_ sky130_fd_sc_hd__a21o_1
X_12820_ _05259_ _05306_ VGND VGND VPWR VPWR _05307_ sky130_fd_sc_hd__xor2_1
XANTENNA__11672__C _06733_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12751_ _05219_ _05229_ VGND VGND VPWR VPWR _05231_ sky130_fd_sc_hd__and2_1
XTAP_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11702_ _04062_ _04067_ VGND VGND VPWR VPWR _04077_ sky130_fd_sc_hd__xnor2_1
XTAP_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_387 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12682_ _05154_ VGND VGND VPWR VPWR _05155_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12784__B _00572_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11633_ _03969_ _03997_ _04000_ VGND VGND VPWR VPWR _04001_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07878__B _06744_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10585__A _02158_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11564_ _01247_ _03914_ _03913_ VGND VGND VPWR VPWR _03925_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_92_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13303_ _05525_ _05595_ _05822_ _05823_ _05824_ VGND VGND VPWR VPWR _05825_ sky130_fd_sc_hd__a311o_4
XFILLER_0_134_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10515_ _02760_ _02764_ VGND VGND VPWR VPWR _02772_ sky130_fd_sc_hd__or2_1
XFILLER_0_107_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11495_ _03846_ _03848_ VGND VGND VPWR VPWR _03849_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07894__A net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13234_ _05575_ _05759_ VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__xnor2_4
XFILLER_0_21_822 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10446_ _02695_ _02472_ _02696_ VGND VGND VPWR VPWR _02698_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_122_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10538__A1 _00293_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10538__B2 _03015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13165_ _05616_ _05463_ _05612_ VGND VGND VPWR VPWR _05686_ sky130_fd_sc_hd__a21oi_2
X_10377_ _03521_ _00734_ VGND VGND VPWR VPWR _02622_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12116_ _04515_ _04516_ VGND VGND VPWR VPWR _04533_ sky130_fd_sc_hd__xnor2_2
X_13096_ _04548_ _04550_ VGND VGND VPWR VPWR _05611_ sky130_fd_sc_hd__nand2_1
XFILLER_0_137_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12047_ _04326_ _04456_ VGND VGND VPWR VPWR _04457_ sky130_fd_sc_hd__xnor2_1
X_13998_ _06556_ _06561_ _06547_ VGND VGND VPWR VPWR _06585_ sky130_fd_sc_hd__o21a_1
XFILLER_0_1_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10479__B _00636_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12949_ _05430_ _05448_ VGND VGND VPWR VPWR _05449_ sky130_fd_sc_hd__or2_1
XFILLER_0_75_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08140_ _06985_ _07082_ VGND VGND VPWR VPWR _00184_ sky130_fd_sc_hd__nand2_1
XFILLER_0_114_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08071_ _01383_ _00114_ VGND VGND VPWR VPWR _00115_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_107 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13715__A1 _02426_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08973_ _00950_ _00951_ VGND VGND VPWR VPWR _01084_ sky130_fd_sc_hd__nand2_1
XANTENNA__09227__C _04015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11476__D _02135_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07924_ _07044_ _07051_ VGND VGND VPWR VPWR _07053_ sky130_fd_sc_hd__or2_1
X_07855_ _06935_ _06983_ VGND VGND VPWR VPWR _06984_ sky130_fd_sc_hd__xor2_2
XFILLER_0_79_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07786_ _01000_ _04378_ VGND VGND VPWR VPWR _06915_ sky130_fd_sc_hd__nand2_1
X_09525_ _01528_ _01687_ VGND VGND VPWR VPWR _01688_ sky130_fd_sc_hd__or2_1
XFILLER_0_94_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07979__A _00541_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09456_ _01610_ _01612_ VGND VGND VPWR VPWR _01614_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_93_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08407_ _00290_ _00327_ VGND VGND VPWR VPWR _00466_ sky130_fd_sc_hd__nor2_1
XANTENNA__11009__A2 _00604_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12206__A1 _00784_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09387_ _01535_ _01537_ VGND VGND VPWR VPWR _01538_ sky130_fd_sc_hd__or2_1
XANTENNA__12206__B2 _00374_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08338_ _00390_ VGND VGND VPWR VPWR _00391_ sky130_fd_sc_hd__buf_6
XFILLER_0_105_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10555__D _01933_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08269_ net145 _00314_ VGND VGND VPWR VPWR _00315_ sky130_fd_sc_hd__nor2_1
XFILLER_0_132_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10300_ _02523_ _02536_ VGND VGND VPWR VPWR _02537_ sky130_fd_sc_hd__xnor2_2
XANTENNA__13706__A1 _01288_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11280_ _03514_ _03533_ VGND VGND VPWR VPWR _03614_ sky130_fd_sc_hd__xnor2_2
XANTENNA__13706__B2 _00416_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09386__A1 _00460_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10231_ _01306_ _00672_ net21 net22 VGND VGND VPWR VPWR _02462_ sky130_fd_sc_hd__and4_1
XFILLER_0_104_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_652 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11667__C _00416_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10571__C _01934_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10162_ _02299_ _02241_ _02384_ VGND VGND VPWR VPWR _02386_ sky130_fd_sc_hd__nand3_1
XFILLER_0_100_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10093_ _02165_ _02166_ _02163_ VGND VGND VPWR VPWR _02310_ sky130_fd_sc_hd__a21o_1
X_13921_ net137 net136 VGND VGND VPWR VPWR _06500_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13852_ _05916_ _05919_ VGND VGND VPWR VPWR _06424_ sky130_fd_sc_hd__nor2_1
XFILLER_0_69_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12803_ _05286_ _05287_ VGND VGND VPWR VPWR _05288_ sky130_fd_sc_hd__or2b_1
X_13783_ _06346_ _06347_ VGND VGND VPWR VPWR _06348_ sky130_fd_sc_hd__or2b_1
X_10995_ _02247_ _02190_ _03299_ VGND VGND VPWR VPWR _03300_ sky130_fd_sc_hd__and3_1
XFILLER_0_85_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12734_ _05182_ _05208_ _05209_ _05210_ _05211_ VGND VGND VPWR VPWR _05212_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_32_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12665_ _04724_ _05135_ VGND VGND VPWR VPWR _05136_ sky130_fd_sc_hd__or2_2
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11616_ _03973_ _03981_ VGND VGND VPWR VPWR _03983_ sky130_fd_sc_hd__or2b_1
XFILLER_0_53_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09074__B1 net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12596_ _00745_ _01059_ VGND VGND VPWR VPWR _05061_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07120__C _00672_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11547_ _06965_ _06966_ _02119_ _02120_ VGND VGND VPWR VPWR _03907_ sky130_fd_sc_hd__nand4_1
XFILLER_0_123_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output98_A net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11478_ _03819_ _03821_ VGND VGND VPWR VPWR _03831_ sky130_fd_sc_hd__xnor2_1
X_13217_ _05655_ _05659_ _05662_ VGND VGND VPWR VPWR _05744_ sky130_fd_sc_hd__or3_1
X_10429_ _02677_ _02678_ VGND VGND VPWR VPWR _02679_ sky130_fd_sc_hd__nand2_1
XANTENNA__11773__A1_N _01996_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14197_ _06621_ _06644_ _06697_ VGND VGND VPWR VPWR _06791_ sky130_fd_sc_hd__or3_2
XFILLER_0_122_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13148_ _05649_ _05651_ VGND VGND VPWR VPWR _05668_ sky130_fd_sc_hd__xor2_2
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11296__D _02737_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13079_ _05548_ _05561_ VGND VGND VPWR VPWR _05592_ sky130_fd_sc_hd__or2b_2
XFILLER_0_79_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07640_ _05709_ _05977_ VGND VGND VPWR VPWR _06373_ sky130_fd_sc_hd__or2b_1
X_07571_ _05621_ _05544_ VGND VGND VPWR VPWR _05632_ sky130_fd_sc_hd__and2b_1
XFILLER_0_88_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09310_ _01450_ _01452_ VGND VGND VPWR VPWR _01453_ sky130_fd_sc_hd__xor2_1
XFILLER_0_48_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09241_ _01366_ _01081_ _01377_ VGND VGND VPWR VPWR _01378_ sky130_fd_sc_hd__o21a_1
XFILLER_0_146_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09460__A2_N _03894_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08407__B _00327_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09172_ _03521_ _00486_ _03707_ _03740_ VGND VGND VPWR VPWR _01302_ sky130_fd_sc_hd__nand4_4
XFILLER_0_56_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_418 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08123_ _00069_ _00165_ VGND VGND VPWR VPWR _00167_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10953__A _00298_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10080__D1 _01486_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08054_ _00000_ _00097_ VGND VGND VPWR VPWR _00098_ sky130_fd_sc_hd__nor2_1
XFILLER_0_113_142 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13686__D _02731_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12590__D _02857_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08956_ _00460_ VGND VGND VPWR VPWR _01066_ sky130_fd_sc_hd__buf_4
X_07907_ _07005_ _07035_ VGND VGND VPWR VPWR _07036_ sky130_fd_sc_hd__xor2_2
X_08887_ _00251_ _00712_ _00985_ _00986_ _00990_ VGND VGND VPWR VPWR _00991_ sky130_fd_sc_hd__a311o_4
XANTENNA__09540__A1 _05192_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07838_ _01383_ _01350_ _06965_ _06966_ VGND VGND VPWR VPWR _06967_ sky130_fd_sc_hd__and4_1
XFILLER_0_98_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11008__B _01505_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07769_ _06723_ _06896_ _06894_ VGND VGND VPWR VPWR _06898_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_39_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09508_ _01668_ _01669_ VGND VGND VPWR VPWR _01670_ sky130_fd_sc_hd__xnor2_1
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10780_ _06637_ _02720_ _03055_ _03054_ VGND VGND VPWR VPWR _03064_ sky130_fd_sc_hd__a31o_1
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07502__A net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09439_ _01582_ _01594_ VGND VGND VPWR VPWR _01595_ sky130_fd_sc_hd__xnor2_1
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12450_ _04824_ _04899_ VGND VGND VPWR VPWR _04900_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11401_ _03743_ _03745_ VGND VGND VPWR VPWR _03746_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_90_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10863__A _05566_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12381_ _04811_ _04821_ _04823_ VGND VGND VPWR VPWR _04824_ sky130_fd_sc_hd__a21oi_1
X_14120_ _06099_ _06656_ _06675_ VGND VGND VPWR VPWR _06717_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_62_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11332_ _03660_ _03670_ VGND VGND VPWR VPWR _03671_ sky130_fd_sc_hd__xnor2_2
XANTENNA__09429__A _01211_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10582__B _01413_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14051_ _06636_ _06642_ VGND VGND VPWR VPWR _06643_ sky130_fd_sc_hd__or2_2
X_11263_ _03032_ _03594_ VGND VGND VPWR VPWR _03595_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08052__B _00095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13002_ _05505_ _05506_ VGND VGND VPWR VPWR _05507_ sky130_fd_sc_hd__and2b_1
X_10214_ _02440_ _02441_ VGND VGND VPWR VPWR _02443_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11194_ _03221_ _03239_ _03241_ VGND VGND VPWR VPWR _03519_ sky130_fd_sc_hd__a21oi_1
X_10145_ _05027_ _04048_ _02365_ _02366_ VGND VGND VPWR VPWR _02367_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_27_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10076_ _02263_ _02266_ _02289_ VGND VGND VPWR VPWR _02292_ sky130_fd_sc_hd__a21o_1
XFILLER_0_89_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12302__B _00575_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13904_ _06433_ _06480_ VGND VGND VPWR VPWR _06481_ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13835_ _06397_ _06402_ _06404_ VGND VGND VPWR VPWR _06405_ sky130_fd_sc_hd__o21ai_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13766_ _06323_ _06327_ _06314_ VGND VGND VPWR VPWR _06330_ sky130_fd_sc_hd__a21oi_1
X_10978_ _03280_ _03281_ VGND VGND VPWR VPWR _03282_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12717_ _05174_ _05176_ VGND VGND VPWR VPWR _05194_ sky130_fd_sc_hd__xor2_2
XFILLER_0_73_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13697_ _00416_ _01288_ _02725_ _02730_ VGND VGND VPWR VPWR _06254_ sky130_fd_sc_hd__and4_1
XFILLER_0_128_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12648_ _05090_ _05117_ VGND VGND VPWR VPWR _05118_ sky130_fd_sc_hd__xor2_2
XFILLER_0_72_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12579_ _00393_ _02758_ _02720_ _00390_ VGND VGND VPWR VPWR _05042_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10601__B1 _02158_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08810_ _00300_ net15 _00732_ _00731_ VGND VGND VPWR VPWR _00906_ sky130_fd_sc_hd__a31o_1
XFILLER_0_110_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09790_ _01977_ _01978_ VGND VGND VPWR VPWR _01979_ sky130_fd_sc_hd__and2b_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08741_ _00543_ _00656_ _00829_ VGND VGND VPWR VPWR _00831_ sky130_fd_sc_hd__a21oi_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09505__C _01508_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08672_ _03894_ VGND VGND VPWR VPWR _00755_ sky130_fd_sc_hd__buf_4
XFILLER_0_84_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07623_ _02007_ _05588_ _05827_ _05818_ VGND VGND VPWR VPWR _06186_ sky130_fd_sc_hd__a31o_1
XFILLER_0_88_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07554_ _01044_ VGND VGND VPWR VPWR _05445_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_76_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07485_ net33 _04455_ VGND VGND VPWR VPWR _04686_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09224_ _01355_ _01358_ VGND VGND VPWR VPWR _01359_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_75_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09155_ _01269_ _01282_ VGND VGND VPWR VPWR _01283_ sky130_fd_sc_hd__xor2_1
XANTENNA__13697__C _02725_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09894__D _02088_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08106_ _00148_ _00149_ VGND VGND VPWR VPWR _00150_ sky130_fd_sc_hd__or2_1
X_09086_ _03850_ _01394_ _00730_ net15 VGND VGND VPWR VPWR _01209_ sky130_fd_sc_hd__and4_1
XFILLER_0_102_602 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08037_ _00080_ VGND VGND VPWR VPWR _00081_ sky130_fd_sc_hd__buf_6
XFILLER_0_4_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08564__A2 _00636_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09988_ _02186_ _02194_ VGND VGND VPWR VPWR _02196_ sky130_fd_sc_hd__nor2_1
XANTENNA__07772__B1 net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08939_ _00991_ _01047_ VGND VGND VPWR VPWR _01048_ sky130_fd_sc_hd__xor2_2
X_11950_ _04271_ _04280_ _04278_ VGND VGND VPWR VPWR _04350_ sky130_fd_sc_hd__a21oi_1
X_10901_ _03194_ _03196_ VGND VGND VPWR VPWR _03197_ sky130_fd_sc_hd__nand2_1
XANTENNA__11961__B _03678_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11881_ _04051_ _04087_ _04089_ _04273_ VGND VGND VPWR VPWR _04274_ sky130_fd_sc_hd__a211o_1
X_13620_ _06118_ _06119_ _06130_ _06168_ VGND VGND VPWR VPWR _06169_ sky130_fd_sc_hd__or4_1
X_10832_ _01339_ net54 VGND VGND VPWR VPWR _03121_ sky130_fd_sc_hd__nand2_1
XANTENNA__08328__A _00379_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13551_ _06018_ _04013_ _06034_ VGND VGND VPWR VPWR _06093_ sky130_fd_sc_hd__and3_1
XFILLER_0_13_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10763_ _03029_ _03042_ _03044_ VGND VGND VPWR VPWR _03045_ sky130_fd_sc_hd__o21a_1
XFILLER_0_82_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07589__D _00650_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08047__B _00377_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12502_ _04048_ _03894_ _04955_ _04956_ VGND VGND VPWR VPWR _04957_ sky130_fd_sc_hd__a31o_1
XFILLER_0_81_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13482_ _06013_ _06015_ _06016_ VGND VGND VPWR VPWR _06017_ sky130_fd_sc_hd__or3b_1
XFILLER_0_125_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10694_ _02964_ _02961_ VGND VGND VPWR VPWR _02969_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11689__A _06819_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12433_ _04879_ _04880_ VGND VGND VPWR VPWR _04881_ sky130_fd_sc_hd__and2_1
XANTENNA__10593__A _02857_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09159__A _00575_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12364_ _00741_ _00457_ VGND VGND VPWR VPWR _04805_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14103_ _06684_ _06690_ VGND VGND VPWR VPWR _06698_ sky130_fd_sc_hd__or2_1
XFILLER_0_50_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11315_ _03643_ _03650_ VGND VGND VPWR VPWR _03652_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12295_ _02188_ _02427_ _02190_ _02088_ VGND VGND VPWR VPWR _04729_ sky130_fd_sc_hd__and4_1
XFILLER_0_120_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14034_ net133 VGND VGND VPWR VPWR _06624_ sky130_fd_sc_hd__inv_2
XANTENNA__08004__A1 _01044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11246_ _03574_ _03562_ _03567_ VGND VGND VPWR VPWR _03577_ sky130_fd_sc_hd__nor3_1
XFILLER_0_129_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11177_ _03386_ _03402_ _03441_ VGND VGND VPWR VPWR _03501_ sky130_fd_sc_hd__and3_1
XANTENNA__09606__B _01600_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10362__A2 _03894_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10128_ _02222_ _02223_ _02225_ _02348_ _02231_ VGND VGND VPWR VPWR _02349_ sky130_fd_sc_hd__a32o_2
X_10059_ _02052_ _02273_ VGND VGND VPWR VPWR _02274_ sky130_fd_sc_hd__xor2_4
XANTENNA__09504__B2 _02116_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13818_ _01400_ _02187_ _03686_ VGND VGND VPWR VPWR _06387_ sky130_fd_sc_hd__and3_1
XFILLER_0_147_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07142__A net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13749_ _06292_ _06309_ _06310_ VGND VGND VPWR VPWR _06311_ sky130_fd_sc_hd__and3_1
XFILLER_0_45_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07270_ _00453_ _02280_ _02313_ VGND VGND VPWR VPWR _02324_ sky130_fd_sc_hd__and3_1
XFILLER_0_85_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13798__B _02190_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_850 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_552 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_782 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12207__B _03682_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09911_ _01978_ _02110_ VGND VGND VPWR VPWR _02111_ sky130_fd_sc_hd__nand2_1
XFILLER_0_111_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10950__B _04906_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09842_ _01825_ _01827_ _02034_ _02035_ VGND VGND VPWR VPWR _02036_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_95_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07962__D _06885_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09773_ net20 VGND VGND VPWR VPWR _01960_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__09235__C _01368_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08724_ _00809_ _00811_ VGND VGND VPWR VPWR _00812_ sky130_fd_sc_hd__or2_1
XTAP_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12666__B1_N _05136_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12877__B _02119_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08655_ _00733_ _00735_ VGND VGND VPWR VPWR _00736_ sky130_fd_sc_hd__xnor2_1
XTAP_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07606_ net191 net192 VGND VGND VPWR VPWR _05999_ sky130_fd_sc_hd__nand2_2
XTAP_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08586_ _00659_ _00660_ VGND VGND VPWR VPWR _00662_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07537_ _04587_ _05247_ _04565_ VGND VGND VPWR VPWR _05258_ sky130_fd_sc_hd__a21o_1
XANTENNA__12893__A _00783_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07468_ _03850_ _01394_ _04378_ _04455_ VGND VGND VPWR VPWR _04499_ sky130_fd_sc_hd__nand4_2
XFILLER_0_9_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09207_ _01144_ _01330_ _01340_ VGND VGND VPWR VPWR _01341_ sky130_fd_sc_hd__and3_1
XFILLER_0_32_500 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07399_ _03729_ VGND VGND VPWR VPWR _03740_ sky130_fd_sc_hd__buf_4
XFILLER_0_106_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09138_ _01263_ _01264_ VGND VGND VPWR VPWR _01265_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09069_ _00913_ _00933_ VGND VGND VPWR VPWR _01190_ sky130_fd_sc_hd__nand2_1
XFILLER_0_130_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09129__D _01254_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11100_ _03277_ _03415_ VGND VGND VPWR VPWR _03416_ sky130_fd_sc_hd__nor2_1
X_12080_ _02246_ _02426_ _04330_ VGND VGND VPWR VPWR _04493_ sky130_fd_sc_hd__and3_1
XFILLER_0_102_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11031_ net7 _00782_ _00778_ _05027_ VGND VGND VPWR VPWR _03340_ sky130_fd_sc_hd__a22oi_1
XANTENNA__11541__A1 _06873_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11541__B2 _06874_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11557__A1_N _03521_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12982_ _05476_ _05484_ VGND VGND VPWR VPWR _05485_ sky130_fd_sc_hd__and2_1
XFILLER_0_99_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11933_ _00113_ _00574_ _04330_ VGND VGND VPWR VPWR _04331_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11864_ _04122_ _04141_ _04254_ VGND VGND VPWR VPWR _04255_ sky130_fd_sc_hd__a21o_1
XANTENNA__08058__A _00628_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13603_ _06138_ _06147_ _06148_ _06149_ VGND VGND VPWR VPWR _06150_ sky130_fd_sc_hd__nor4_1
X_10815_ _06937_ _02735_ VGND VGND VPWR VPWR _03102_ sky130_fd_sc_hd__nand2_1
XANTENNA__13597__A2 _01249_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11795_ _01361_ _00159_ _02459_ _02673_ VGND VGND VPWR VPWR _04179_ sky130_fd_sc_hd__nand4_1
XFILLER_0_55_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13534_ _02766_ VGND VGND VPWR VPWR _06074_ sky130_fd_sc_hd__buf_2
XFILLER_0_39_187 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10746_ _03008_ _03010_ VGND VGND VPWR VPWR _03027_ sky130_fd_sc_hd__xor2_1
XFILLER_0_94_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13465_ _05996_ _05997_ VGND VGND VPWR VPWR _05998_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10677_ _05181_ _01411_ VGND VGND VPWR VPWR _02951_ sky130_fd_sc_hd__nand2_1
X_12416_ _00378_ _01586_ VGND VGND VPWR VPWR _04863_ sky130_fd_sc_hd__nand2_2
XFILLER_0_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13396_ _05921_ _05922_ VGND VGND VPWR VPWR _05924_ sky130_fd_sc_hd__or2_1
XFILLER_0_51_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12347_ _04783_ _04786_ VGND VGND VPWR VPWR _04787_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_output80_A net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11866__B _00258_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12278_ _04701_ _04710_ VGND VGND VPWR VPWR _04711_ sky130_fd_sc_hd__and2b_1
XFILLER_0_121_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14017_ _06599_ _06602_ VGND VGND VPWR VPWR _06606_ sky130_fd_sc_hd__or2b_1
X_11229_ _03434_ _03436_ _03430_ VGND VGND VPWR VPWR _03558_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07137__A net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11882__A _00262_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08440_ _02018_ _00158_ _00501_ VGND VGND VPWR VPWR _00502_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11106__B _01066_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08371_ _01744_ net11 _00422_ _00424_ VGND VGND VPWR VPWR _00426_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__13588__A2 _03783_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07303__C _00573_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07322_ _02445_ _02883_ VGND VGND VPWR VPWR _02894_ sky130_fd_sc_hd__nand2_2
XFILLER_0_18_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_95 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07253_ _02127_ VGND VGND VPWR VPWR _02138_ sky130_fd_sc_hd__buf_4
XFILLER_0_6_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07184_ _01372_ VGND VGND VPWR VPWR _01383_ sky130_fd_sc_hd__buf_6
XFILLER_0_131_516 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11771__A1 _05445_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11771__B2 _05467_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11776__B _05478_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10680__B _02982_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13512__A2 _02736_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09825_ _03510_ net11 VGND VGND VPWR VPWR _02017_ sky130_fd_sc_hd__nand2_1
XANTENNA__12888__A _00379_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09756_ _01889_ _01940_ VGND VGND VPWR VPWR _01942_ sky130_fd_sc_hd__xnor2_1
X_08707_ _00791_ _00793_ VGND VGND VPWR VPWR _00794_ sky130_fd_sc_hd__and2b_1
XFILLER_0_69_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09687_ _01862_ _01863_ VGND VGND VPWR VPWR _01866_ sky130_fd_sc_hd__and2_1
XTAP_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08638_ _00439_ _00560_ _00559_ VGND VGND VPWR VPWR _00719_ sky130_fd_sc_hd__a21oi_2
XTAP_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10201__A _06626_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08569_ _03543_ _00294_ _00533_ _00532_ VGND VGND VPWR VPWR _00643_ sky130_fd_sc_hd__a31o_1
XFILLER_0_77_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10600_ _04862_ _04873_ _01410_ _02158_ VGND VGND VPWR VPWR _02866_ sky130_fd_sc_hd__and4_1
X_11580_ _03893_ _03941_ _03942_ VGND VGND VPWR VPWR _03943_ sky130_fd_sc_hd__or3_1
XFILLER_0_119_362 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_682 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10855__B _02855_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10531_ _02754_ _02756_ _02789_ VGND VGND VPWR VPWR _02790_ sky130_fd_sc_hd__a21o_1
XFILLER_0_24_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13250_ _01647_ _01648_ _05774_ _05775_ VGND VGND VPWR VPWR _05776_ sky130_fd_sc_hd__a211o_4
X_10462_ _02052_ _02273_ _02279_ VGND VGND VPWR VPWR _02715_ sky130_fd_sc_hd__a21o_1
XFILLER_0_17_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12201_ _03667_ _04625_ VGND VGND VPWR VPWR _04626_ sky130_fd_sc_hd__xor2_2
XANTENNA__11211__B1 _02582_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13181_ _04551_ _05703_ VGND VGND VPWR VPWR _05704_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_20_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10393_ _02635_ _02636_ _02634_ VGND VGND VPWR VPWR _02639_ sky130_fd_sc_hd__and3_1
XANTENNA__07966__B1 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12132_ _04523_ _04528_ _04549_ VGND VGND VPWR VPWR _04550_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_32_396 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07883__C net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12063_ _04461_ _04464_ VGND VGND VPWR VPWR _04474_ sky130_fd_sc_hd__or2_1
XANTENNA__12711__B1 _01415_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11014_ _03316_ _03319_ _03320_ VGND VGND VPWR VPWR _03321_ sky130_fd_sc_hd__and3_1
XANTENNA__12798__A _00916_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09172__A _03521_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12965_ _05465_ _03623_ VGND VGND VPWR VPWR _05466_ sky130_fd_sc_hd__xor2_2
XFILLER_0_99_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11916_ _04306_ _04311_ VGND VGND VPWR VPWR _04313_ sky130_fd_sc_hd__nor2_1
XANTENNA__07404__B _01470_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12896_ _05388_ _05389_ VGND VGND VPWR VPWR _05391_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_74_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11847_ _04236_ VGND VGND VPWR VPWR _04237_ sky130_fd_sc_hd__inv_2
XTAP_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_580 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11778_ _04152_ _04154_ _04159_ _04160_ VGND VGND VPWR VPWR _04161_ sky130_fd_sc_hd__o211a_1
XFILLER_0_138_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13517_ _05992_ _06007_ _06005_ VGND VGND VPWR VPWR _06056_ sky130_fd_sc_hd__a21oi_1
X_10729_ _02835_ _03007_ VGND VGND VPWR VPWR _03008_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10484__C _02736_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13448_ _01252_ _02736_ _02731_ _01182_ VGND VGND VPWR VPWR _05980_ sky130_fd_sc_hd__a22o_1
XFILLER_0_140_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10781__A _06937_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13379_ _05903_ _05904_ VGND VGND VPWR VPWR _05905_ sky130_fd_sc_hd__nand2_1
XANTENNA__07957__B1 _03015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08889__C _04906_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08251__A _06428_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07940_ _07055_ _07068_ VGND VGND VPWR VPWR _07069_ sky130_fd_sc_hd__nor2_1
X_07871_ _06998_ _06999_ VGND VGND VPWR VPWR _07000_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10005__B _04598_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09610_ _02280_ _01780_ _01781_ VGND VGND VPWR VPWR _01782_ sky130_fd_sc_hd__and3_1
XANTENNA__12501__A _04026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09541_ _04598_ net40 VGND VGND VPWR VPWR _01706_ sky130_fd_sc_hd__nand2_1
XFILLER_0_116_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09472_ _01627_ _01628_ _01629_ _01630_ VGND VGND VPWR VPWR _01631_ sky130_fd_sc_hd__o211a_1
XFILLER_0_78_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08423_ _00280_ _00482_ VGND VGND VPWR VPWR _00483_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10956__A _04895_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_660 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08354_ _00395_ _00407_ VGND VGND VPWR VPWR _00408_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08437__A1 _05456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_742 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07305_ _02686_ _02697_ VGND VGND VPWR VPWR _02708_ sky130_fd_sc_hd__and2b_1
XANTENNA__07330__A _02971_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08285_ _00330_ _00331_ VGND VGND VPWR VPWR _00332_ sky130_fd_sc_hd__or2b_1
XFILLER_0_74_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07236_ _00694_ _01941_ VGND VGND VPWR VPWR _01952_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07167_ net58 VGND VGND VPWR VPWR _01197_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__14163__A _02742_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07098_ _00431_ VGND VGND VPWR VPWR _00442_ sky130_fd_sc_hd__buf_6
XFILLER_0_112_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09808_ _01791_ _01794_ _01790_ VGND VGND VPWR VPWR _01999_ sky130_fd_sc_hd__o21a_1
XANTENNA__09704__B _00459_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12411__A _00378_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07505__A _04895_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09739_ _04169_ _01076_ _01545_ net52 VGND VGND VPWR VPWR _01923_ sky130_fd_sc_hd__and4_1
XANTENNA__11672__D net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12750_ _05219_ _05229_ VGND VGND VPWR VPWR _05230_ sky130_fd_sc_hd__nor2_1
XTAP_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11701_ _02625_ _02624_ VGND VGND VPWR VPWR _04076_ sky130_fd_sc_hd__or2b_1
XTAP_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12681_ _05145_ _05150_ _05152_ _05153_ VGND VGND VPWR VPWR _05154_ sky130_fd_sc_hd__o211a_1
XTAP_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12784__C _01411_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11632_ _03998_ _03999_ VGND VGND VPWR VPWR _04000_ sky130_fd_sc_hd__nand2_1
XTAP_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_107 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08336__A _03707_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07240__A _01000_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11563_ _03917_ _03922_ _03923_ VGND VGND VPWR VPWR _03924_ sky130_fd_sc_hd__nor3_1
XFILLER_0_65_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_639 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13302_ _05603_ _05822_ VGND VGND VPWR VPWR _05824_ sky130_fd_sc_hd__and2_1
XFILLER_0_107_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10514_ _02247_ _02765_ VGND VGND VPWR VPWR _02771_ sky130_fd_sc_hd__nand2_1
XFILLER_0_107_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11494_ _03838_ _03847_ VGND VGND VPWR VPWR _03848_ sky130_fd_sc_hd__or2_1
XFILLER_0_134_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13233_ _02278_ _05756_ _05758_ VGND VGND VPWR VPWR _05759_ sky130_fd_sc_hd__a21oi_2
XANTENNA__07894__B net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10445_ _02424_ _02437_ VGND VGND VPWR VPWR _02696_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10538__A2 _02725_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_480 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13164_ _03493_ _05684_ VGND VGND VPWR VPWR _05685_ sky130_fd_sc_hd__xnor2_4
XANTENNA__08071__A _01383_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10376_ _00413_ _02618_ _02619_ VGND VGND VPWR VPWR _02621_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_103_571 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12115_ _04519_ _04530_ VGND VGND VPWR VPWR _04531_ sky130_fd_sc_hd__xor2_4
X_13095_ _03956_ _04025_ _04545_ VGND VGND VPWR VPWR _05609_ sky130_fd_sc_hd__nor3b_1
X_12046_ _04253_ _04322_ VGND VGND VPWR VPWR _04456_ sky130_fd_sc_hd__xor2_1
XFILLER_0_137_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13997_ _06583_ VGND VGND VPWR VPWR _06584_ sky130_fd_sc_hd__inv_2
XANTENNA__10479__C _02726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12948_ _05435_ _05447_ VGND VGND VPWR VPWR _05448_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13660__A1 _01415_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09864__B1 _00393_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13660__B2 _01108_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11671__B1 _03762_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12879_ _05369_ _05370_ _05371_ VGND VGND VPWR VPWR _05372_ sky130_fd_sc_hd__a21oi_1
XTAP_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__07150__A _00442_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_786 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08070_ _00101_ VGND VGND VPWR VPWR _00114_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_114_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13715__A2 _02759_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11400__A _00003_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12215__B _03750_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08972_ _01081_ _01082_ VGND VGND VPWR VPWR _01083_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07923_ _07044_ _07051_ VGND VGND VPWR VPWR _07052_ sky130_fd_sc_hd__and2_1
XFILLER_0_39_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07854_ _06981_ _06982_ VGND VGND VPWR VPWR _06983_ sky130_fd_sc_hd__nand2_2
XANTENNA__13046__B _05554_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07785_ _06912_ _06913_ VGND VGND VPWR VPWR _06914_ sky130_fd_sc_hd__and2b_1
XFILLER_0_78_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09524_ _01501_ _01526_ _01538_ VGND VGND VPWR VPWR _01687_ sky130_fd_sc_hd__o21a_1
X_09455_ _01187_ _01227_ _01297_ _01611_ VGND VGND VPWR VPWR _01612_ sky130_fd_sc_hd__a31o_4
XANTENNA__07979__B _02719_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10686__A _05181_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08406_ _00254_ _00328_ VGND VGND VPWR VPWR _00465_ sky130_fd_sc_hd__nor2_1
XFILLER_0_143_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09386_ _00460_ _01399_ _01534_ VGND VGND VPWR VPWR _01537_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12206__A2 _01953_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08337_ _00389_ VGND VGND VPWR VPWR _00390_ sky130_fd_sc_hd__buf_4
XFILLER_0_47_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_611 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08268_ _00306_ _00307_ _00309_ _00312_ VGND VGND VPWR VPWR _00314_ sky130_fd_sc_hd__o22a_1
XFILLER_0_117_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07219_ _01733_ _01755_ VGND VGND VPWR VPWR _01766_ sky130_fd_sc_hd__nand2_1
XANTENNA__13706__A2 _02720_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08199_ _00190_ _00191_ _00201_ VGND VGND VPWR VPWR _00243_ sky130_fd_sc_hd__and3_1
XFILLER_0_30_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10230_ _02460_ VGND VGND VPWR VPWR _02461_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11667__D _01288_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10571__D _02169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10161_ _02299_ _02241_ _02384_ VGND VGND VPWR VPWR _02385_ sky130_fd_sc_hd__a21o_1
XANTENNA__09715__A _06483_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10092_ _02303_ _02308_ VGND VGND VPWR VPWR _02309_ sky130_fd_sc_hd__xor2_2
X_13920_ _06496_ _06498_ VGND VGND VPWR VPWR _06499_ sky130_fd_sc_hd__nand2_1
X_13851_ _05904_ _06420_ _06422_ VGND VGND VPWR VPWR _06423_ sky130_fd_sc_hd__and3_1
X_12802_ _05106_ _05285_ VGND VGND VPWR VPWR _05287_ sky130_fd_sc_hd__nand2_1
X_13782_ _05884_ _05889_ _05885_ VGND VGND VPWR VPWR _06347_ sky130_fd_sc_hd__o21ai_1
X_10994_ _01473_ _02188_ VGND VGND VPWR VPWR _03299_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12733_ _05173_ _05180_ VGND VGND VPWR VPWR _05211_ sky130_fd_sc_hd__or2_1
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12664_ _04721_ _04723_ VGND VGND VPWR VPWR _05135_ sky130_fd_sc_hd__and2_1
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11615_ _03977_ _03979_ _03980_ VGND VGND VPWR VPWR _03981_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_5_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09074__A1 _05445_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09074__B2 _05731_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12595_ _05052_ _05058_ VGND VGND VPWR VPWR _05059_ sky130_fd_sc_hd__xor2_2
XFILLER_0_37_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11546_ _03532_ _02120_ _03900_ _03899_ VGND VGND VPWR VPWR _03906_ sky130_fd_sc_hd__a31o_1
XFILLER_0_25_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07120__D _00300_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11477_ _03827_ _03829_ VGND VGND VPWR VPWR _03830_ sky130_fd_sc_hd__and2_1
XFILLER_0_80_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13216_ _05713_ _05737_ _05741_ VGND VGND VPWR VPWR _05743_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_123_699 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10428_ _02671_ _02676_ VGND VGND VPWR VPWR _02678_ sky130_fd_sc_hd__or2_1
X_14196_ _06621_ _06778_ VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__xnor2_4
XFILLER_0_21_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13147_ _05664_ _05659_ _05666_ _05658_ VGND VGND VPWR VPWR _05667_ sky130_fd_sc_hd__a22o_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10359_ _03696_ _02600_ _02601_ VGND VGND VPWR VPWR _02602_ sky130_fd_sc_hd__a21bo_1
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13078_ _05590_ _05578_ _05574_ VGND VGND VPWR VPWR _05591_ sky130_fd_sc_hd__a21o_1
XFILLER_0_57_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12029_ _04365_ _04435_ VGND VGND VPWR VPWR _04437_ sky130_fd_sc_hd__nor2_1
X_07570_ _05555_ _05610_ VGND VGND VPWR VPWR _05621_ sky130_fd_sc_hd__xor2_2
XFILLER_0_73_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09360__A _01507_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09240_ _01375_ _01376_ VGND VGND VPWR VPWR _01377_ sky130_fd_sc_hd__nor2_1
XFILLER_0_146_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09171_ _03554_ _00391_ _00393_ _00519_ VGND VGND VPWR VPWR _01301_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08122_ _00069_ _00165_ VGND VGND VPWR VPWR _00166_ sky130_fd_sc_hd__and2_1
XANTENNA__08704__A _00442_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10953__B _00608_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08053_ _00093_ _00096_ VGND VGND VPWR VPWR _00097_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12226__A _01518_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09535__A _00355_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08955_ _00981_ _00983_ _01063_ VGND VGND VPWR VPWR _01064_ sky130_fd_sc_hd__a21o_1
X_07906_ _07033_ _07034_ VGND VGND VPWR VPWR _07035_ sky130_fd_sc_hd__or2b_1
X_08886_ _00881_ _00987_ _00988_ VGND VGND VPWR VPWR _00990_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10135__B1 _01368_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09540__A2 net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07837_ _06875_ VGND VGND VPWR VPWR _06966_ sky130_fd_sc_hd__clkbuf_4
X_07768_ _06723_ _06894_ _06896_ VGND VGND VPWR VPWR _06897_ sky130_fd_sc_hd__and3_1
XFILLER_0_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09270__A net50 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09507_ _06472_ _00607_ VGND VGND VPWR VPWR _01669_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07699_ _06809_ _06816_ _06826_ VGND VGND VPWR VPWR _06828_ sky130_fd_sc_hd__a21oi_1
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09438_ _01592_ _01593_ VGND VGND VPWR VPWR _01594_ sky130_fd_sc_hd__and2_1
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09369_ _00784_ VGND VGND VPWR VPWR _01518_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_136_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11400_ _00003_ _03744_ VGND VGND VPWR VPWR _03745_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12380_ _04798_ _04822_ VGND VGND VPWR VPWR _04823_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11331_ _03661_ _03658_ VGND VGND VPWR VPWR _03670_ sky130_fd_sc_hd__and2_1
XFILLER_0_132_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14050_ _06641_ VGND VGND VPWR VPWR _06642_ sky130_fd_sc_hd__inv_2
X_11262_ _02980_ _02983_ VGND VGND VPWR VPWR _03594_ sky130_fd_sc_hd__and2_1
XANTENNA__07586__A1_N _02029_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13001_ _05504_ _05496_ _05502_ VGND VGND VPWR VPWR _05506_ sky130_fd_sc_hd__nand3b_2
XANTENNA__12363__A1 _00755_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10213_ _02440_ _02441_ VGND VGND VPWR VPWR _02442_ sky130_fd_sc_hd__and2_1
XFILLER_0_120_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11193_ _03516_ _03517_ VGND VGND VPWR VPWR _03518_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09445__A _01600_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10144_ _04851_ net4 _04015_ _00780_ VGND VGND VPWR VPWR _02366_ sky130_fd_sc_hd__and4_1
XFILLER_0_100_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10075_ _02263_ _02266_ _02289_ VGND VGND VPWR VPWR _02290_ sky130_fd_sc_hd__and3_1
XANTENNA__12302__C _01664_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13903_ _06416_ _06434_ VGND VGND VPWR VPWR _06480_ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13834_ _06382_ _06403_ VGND VGND VPWR VPWR _06404_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13765_ _06314_ _06323_ _06327_ VGND VGND VPWR VPWR _06328_ sky130_fd_sc_hd__and3_1
XANTENNA__09295__A1 _00898_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10977_ _00143_ _00607_ VGND VGND VPWR VPWR _03281_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12716_ _05183_ _05186_ _05187_ _05189_ _05191_ VGND VGND VPWR VPWR _05193_ sky130_fd_sc_hd__a32oi_4
XFILLER_0_45_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13696_ _06250_ _06251_ VGND VGND VPWR VPWR _06253_ sky130_fd_sc_hd__and2_1
XFILLER_0_26_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12647_ _05099_ _05116_ VGND VGND VPWR VPWR _05117_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_115_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12578_ _05040_ VGND VGND VPWR VPWR _05041_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10601__A1 _04862_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11529_ _03880_ _03882_ VGND VGND VPWR VPWR _03887_ sky130_fd_sc_hd__or2_1
XANTENNA__10601__B2 _04873_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14179_ _06763_ _06766_ VGND VGND VPWR VPWR _06779_ sky130_fd_sc_hd__and2_1
XFILLER_0_68_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08740_ _07004_ _00656_ _00829_ VGND VGND VPWR VPWR _00830_ sky130_fd_sc_hd__and3_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09505__D _01504_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08671_ _00752_ _00753_ VGND VGND VPWR VPWR _00754_ sky130_fd_sc_hd__or2b_1
XFILLER_0_108_62 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07622_ _06076_ _06164_ net183 VGND VGND VPWR VPWR _06175_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_17_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13606__A1 _02856_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07553_ _03136_ _03158_ _03169_ VGND VGND VPWR VPWR _05434_ sky130_fd_sc_hd__and3_1
XFILLER_0_49_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11770__D net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07484_ _04653_ _04664_ VGND VGND VPWR VPWR _04675_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_124_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_818 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09223_ _00991_ _01356_ _01357_ VGND VGND VPWR VPWR _01358_ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_851 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09154_ _01280_ _01281_ VGND VGND VPWR VPWR _01282_ sky130_fd_sc_hd__nor2_1
XANTENNA__13697__D _02730_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08105_ _00045_ _00147_ VGND VGND VPWR VPWR _00149_ sky130_fd_sc_hd__and2_1
XFILLER_0_31_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09085_ _02127_ _00734_ _00902_ _00900_ VGND VGND VPWR VPWR _01207_ sky130_fd_sc_hd__a31o_1
XFILLER_0_102_614 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08036_ _00041_ _00042_ _00078_ _00079_ VGND VGND VPWR VPWR _00080_ sky130_fd_sc_hd__or4_4
XFILLER_0_114_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11795__A _01361_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09987_ _02186_ _02194_ VGND VGND VPWR VPWR _02195_ sky130_fd_sc_hd__and2_1
XANTENNA__07772__A1 _01208_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08938_ _01042_ _01046_ VGND VGND VPWR VPWR _01047_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_99_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08869_ _00969_ _00970_ VGND VGND VPWR VPWR _00971_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10900_ _03164_ _03195_ VGND VGND VPWR VPWR _03196_ sky130_fd_sc_hd__nor2_1
XANTENNA__09712__B _06461_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11880_ _00257_ _00670_ _00915_ _00916_ VGND VGND VPWR VPWR _04273_ sky130_fd_sc_hd__and4_1
XFILLER_0_98_258 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07513__A _00573_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10831_ _03110_ _03109_ VGND VGND VPWR VPWR _03120_ sky130_fd_sc_hd__and2b_1
XFILLER_0_39_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11035__A _00298_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13550_ _06033_ _06039_ _06064_ VGND VGND VPWR VPWR _06092_ sky130_fd_sc_hd__and3_1
XFILLER_0_67_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10762_ _03016_ _03043_ VGND VGND VPWR VPWR _03044_ sky130_fd_sc_hd__nor2_1
XFILLER_0_109_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08047__C _02982_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12501_ _04026_ _00780_ _03685_ _00423_ VGND VGND VPWR VPWR _04956_ sky130_fd_sc_hd__and4_1
XFILLER_0_109_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13481_ _01062_ _01415_ _01958_ _03690_ VGND VGND VPWR VPWR _06016_ sky130_fd_sc_hd__and4_1
XFILLER_0_109_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10693_ _02966_ _02967_ VGND VGND VPWR VPWR _02968_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12432_ _04777_ _04878_ VGND VGND VPWR VPWR _04880_ sky130_fd_sc_hd__or2_1
XFILLER_0_124_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11689__B _06821_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08344__A _00354_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12363_ _00755_ _00457_ _04802_ _04803_ VGND VGND VPWR VPWR _04804_ sky130_fd_sc_hd__a31o_1
XFILLER_0_22_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10595__B1 _02857_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14102_ _05825_ _06695_ _06696_ VGND VGND VPWR VPWR _06697_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_133_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11314_ _03643_ _03650_ VGND VGND VPWR VPWR _03651_ sky130_fd_sc_hd__or2_1
X_12294_ _03414_ _02426_ _04726_ _04727_ VGND VGND VPWR VPWR _04728_ sky130_fd_sc_hd__a31o_1
XFILLER_0_132_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14033_ _06621_ _06622_ VGND VGND VPWR VPWR _06623_ sky130_fd_sc_hd__or2_1
X_11245_ _03562_ _03567_ _03574_ VGND VGND VPWR VPWR _03575_ sky130_fd_sc_hd__o21a_1
XANTENNA__08004__A2 _04367_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11176_ _03189_ _03205_ _03242_ VGND VGND VPWR VPWR _03500_ sky130_fd_sc_hd__and3_1
X_10127_ _02222_ _02227_ VGND VGND VPWR VPWR _02348_ sky130_fd_sc_hd__or2b_1
XANTENNA__09504__A2 _01664_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10058_ _02055_ _02272_ VGND VGND VPWR VPWR _02273_ sky130_fd_sc_hd__xor2_4
XFILLER_0_89_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13817_ _06382_ _06385_ VGND VGND VPWR VPWR _06386_ sky130_fd_sc_hd__and2b_1
XFILLER_0_58_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13748_ _06277_ _06283_ VGND VGND VPWR VPWR _06310_ sky130_fd_sc_hd__xor2_1
XFILLER_0_128_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13679_ _06232_ _06233_ VGND VGND VPWR VPWR _06234_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_564 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08254__A _00158_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12207__C _00379_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_794 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09910_ _00333_ _01955_ _01977_ VGND VGND VPWR VPWR _02110_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10950__C _01508_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07203__B1 _00661_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09841_ _01822_ _01824_ VGND VGND VPWR VPWR _02035_ sky130_fd_sc_hd__nor2_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12315__A2_N _01601_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09772_ _00344_ _01958_ VGND VGND VPWR VPWR _01959_ sky130_fd_sc_hd__nand2_1
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09235__D _00959_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08723_ _00508_ _00144_ _00807_ _00810_ VGND VGND VPWR VPWR _00811_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_21_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08654_ _00311_ _00734_ VGND VGND VPWR VPWR _00735_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07605_ _05709_ _05977_ VGND VGND VPWR VPWR _05988_ sky130_fd_sc_hd__or2_4
XANTENNA__07333__A _03004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13054__B _05554_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08585_ _00653_ _00655_ _00657_ VGND VGND VPWR VPWR _00660_ sky130_fd_sc_hd__and3_1
XTAP_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07536_ _04730_ _04796_ _04807_ VGND VGND VPWR VPWR _05247_ sky130_fd_sc_hd__a21o_1
XFILLER_0_147_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12893__B _00778_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07467_ _00661_ _04455_ _04433_ _04422_ VGND VGND VPWR VPWR _04488_ sky130_fd_sc_hd__a31o_1
XFILLER_0_76_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09206_ _01337_ _01338_ VGND VGND VPWR VPWR _01340_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07398_ _03718_ VGND VGND VPWR VPWR _03729_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_72_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09137_ _01259_ _01261_ _01194_ _01196_ VGND VGND VPWR VPWR _01264_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_32_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09068_ _02456_ _01188_ VGND VGND VPWR VPWR _01189_ sky130_fd_sc_hd__nand2_1
XFILLER_0_130_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_718 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08019_ _00061_ _00062_ VGND VGND VPWR VPWR _00063_ sky130_fd_sc_hd__or2_1
X_11030_ _05027_ net7 _00612_ _00613_ VGND VGND VPWR VPWR _03339_ sky130_fd_sc_hd__and4_1
XANTENNA__07508__A _04928_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12981_ _05480_ _05483_ VGND VGND VPWR VPWR _05484_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11691__C _03510_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11932_ _00114_ _01272_ VGND VGND VPWR VPWR _04330_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08339__A _03740_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__07243__A _00901_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11863_ _04106_ _04121_ VGND VGND VPWR VPWR _04254_ sky130_fd_sc_hd__and2b_1
XFILLER_0_39_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08058__B _00650_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10814_ _03073_ _03100_ VGND VGND VPWR VPWR _03101_ sky130_fd_sc_hd__nor2_1
X_13602_ _01061_ _03783_ _06146_ VGND VGND VPWR VPWR _06149_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11794_ _04172_ _04177_ VGND VGND VPWR VPWR _04178_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13533_ _06071_ _06072_ VGND VGND VPWR VPWR _06073_ sky130_fd_sc_hd__and2_1
XFILLER_0_137_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10745_ _03021_ _03023_ _03024_ VGND VGND VPWR VPWR _03025_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_39_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13464_ _01252_ _05969_ _02735_ _02731_ VGND VGND VPWR VPWR _05997_ sky130_fd_sc_hd__and4_1
XFILLER_0_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10676_ _02941_ _02940_ VGND VGND VPWR VPWR _02950_ sky130_fd_sc_hd__or2b_1
XFILLER_0_51_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_512 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12415_ _04853_ _04852_ VGND VGND VPWR VPWR _04861_ sky130_fd_sc_hd__or2b_2
XFILLER_0_51_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13395_ _05915_ _05920_ VGND VGND VPWR VPWR _05922_ sky130_fd_sc_hd__nor2_1
XFILLER_0_140_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_534 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12346_ _00916_ _01505_ _04784_ VGND VGND VPWR VPWR _04786_ sky130_fd_sc_hd__and3_1
XFILLER_0_11_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12277_ _04705_ _04707_ _04709_ VGND VGND VPWR VPWR _04710_ sky130_fd_sc_hd__a21bo_1
XANTENNA__11866__C _00415_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14016_ _06603_ VGND VGND VPWR VPWR _06605_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_output73_A net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11228_ _03430_ _03434_ _03436_ VGND VGND VPWR VPWR _03557_ sky130_fd_sc_hd__and3_1
XANTENNA__07418__A _00311_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11159_ _03475_ _03480_ VGND VGND VPWR VPWR _03481_ sky130_fd_sc_hd__nand2_2
XANTENNA__11882__B _00263_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08249__A _00095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07153__A net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08370_ _00422_ _00424_ _00672_ net11 VGND VGND VPWR VPWR _00425_ sky130_fd_sc_hd__and4bb_1
XANTENNA__12245__B1 _01248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07303__D net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07321_ _02478_ _02872_ VGND VGND VPWR VPWR _02883_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_45_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_795 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07252_ _00672_ VGND VGND VPWR VPWR _02127_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_26_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07183_ _00891_ VGND VGND VPWR VPWR _01372_ sky130_fd_sc_hd__buf_4
XANTENNA__10019__A _04862_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_720 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11776__C _02117_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09824_ _02013_ _02014_ _02015_ VGND VGND VPWR VPWR _02016_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12888__B _03678_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09755_ _01916_ _01939_ VGND VGND VPWR VPWR _01940_ sky130_fd_sc_hd__xor2_1
X_08706_ _03587_ net46 net47 _00431_ VGND VGND VPWR VPWR _00793_ sky130_fd_sc_hd__a22o_1
X_09686_ _01862_ _01863_ VGND VGND VPWR VPWR _01865_ sky130_fd_sc_hd__nor2_1
XTAP_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08637_ _00598_ _00717_ VGND VGND VPWR VPWR _00718_ sky130_fd_sc_hd__xnor2_2
XTAP_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10201__B _02426_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08568_ _00531_ _00536_ VGND VGND VPWR VPWR _00642_ sky130_fd_sc_hd__nand2_1
XTAP_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07519_ _04884_ _05049_ VGND VGND VPWR VPWR _05060_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08499_ _00565_ _00566_ VGND VGND VPWR VPWR _00567_ sky130_fd_sc_hd__nor2_2
XFILLER_0_37_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12409__A _04059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10530_ _02757_ _02788_ VGND VGND VPWR VPWR _02789_ sky130_fd_sc_hd__nor2_1
XFILLER_0_107_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10461_ _02274_ _02491_ VGND VGND VPWR VPWR _02714_ sky130_fd_sc_hd__and2_1
XFILLER_0_122_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12200_ _03053_ _03673_ _04624_ VGND VGND VPWR VPWR _04625_ sky130_fd_sc_hd__or3b_1
X_13180_ _05482_ _05701_ _04537_ _05702_ _04591_ VGND VGND VPWR VPWR _05703_ sky130_fd_sc_hd__o311a_2
X_10392_ _02634_ _02637_ VGND VGND VPWR VPWR _02638_ sky130_fd_sc_hd__and2b_1
XFILLER_0_60_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07966__A1 _01076_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12131_ _04523_ _04528_ _04522_ VGND VGND VPWR VPWR _04549_ sky130_fd_sc_hd__a21o_1
XANTENNA__07966__B2 _01120_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12144__A _00530_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07883__D net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12062_ _04467_ _04472_ VGND VGND VPWR VPWR _04473_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11013_ _03308_ _03311_ VGND VGND VPWR VPWR _03320_ sky130_fd_sc_hd__xor2_1
XANTENNA__12711__A1 _00393_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12711__B2 _00391_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12798__B _01933_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09172__B _00486_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12964_ _03536_ _03616_ _03621_ VGND VGND VPWR VPWR _05465_ sky130_fd_sc_hd__or3_2
XANTENNA__08069__A _00112_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11915_ _04308_ _04310_ VGND VGND VPWR VPWR _04311_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output111_A net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07404__C _03685_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12895_ _00375_ _02673_ VGND VGND VPWR VPWR _05389_ sky130_fd_sc_hd__nand2_1
XANTENNA__09891__A1 _03070_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11846_ _02456_ _01955_ VGND VGND VPWR VPWR _04236_ sky130_fd_sc_hd__nand2_2
XFILLER_0_51_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_592 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11777_ _05456_ _02117_ _01960_ _05478_ VGND VGND VPWR VPWR _04160_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13516_ _06002_ _06053_ VGND VGND VPWR VPWR _06055_ sky130_fd_sc_hd__xor2_1
X_10728_ _02833_ _02834_ VGND VGND VPWR VPWR _03007_ sky130_fd_sc_hd__or2_1
XFILLER_0_82_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_106 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10484__D _02737_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10659_ _02924_ _02926_ VGND VGND VPWR VPWR _02931_ sky130_fd_sc_hd__nor2_1
X_13447_ _01182_ _01252_ _02735_ _02731_ VGND VGND VPWR VPWR _05979_ sky130_fd_sc_hd__and4_1
XFILLER_0_140_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13378_ _01664_ _01505_ _03738_ _03744_ VGND VGND VPWR VPWR _05904_ sky130_fd_sc_hd__nand4_1
XANTENNA__08532__A _02105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10781__B _06494_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07957__A1 _03554_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07957__B2 _00519_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08889__D _04928_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12329_ _04765_ _04766_ VGND VGND VPWR VPWR _04767_ sky130_fd_sc_hd__and2b_1
XFILLER_0_121_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08251__B _06450_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10961__B1 _02190_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07148__A _00978_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07870_ _06984_ _06899_ VGND VGND VPWR VPWR _06999_ sky130_fd_sc_hd__xor2_2
XANTENNA__10005__C _00782_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09540_ _05192_ net40 _01494_ _01704_ VGND VGND VPWR VPWR _01705_ sky130_fd_sc_hd__a31o_1
XFILLER_0_78_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09471_ _01359_ _01425_ _01309_ VGND VGND VPWR VPWR _01630_ sky130_fd_sc_hd__a21o_1
X_08422_ _00470_ _00481_ VGND VGND VPWR VPWR _00482_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07893__B1 _06820_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10956__B _04873_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08353_ _00384_ _00386_ VGND VGND VPWR VPWR _00407_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08437__A2 _04895_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12229__A _01518_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_683 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07304_ _00705_ _00639_ _00573_ net29 VGND VGND VPWR VPWR _02697_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08284_ _00377_ _06873_ _06875_ _02993_ VGND VGND VPWR VPWR _00331_ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07235_ _00617_ _00683_ VGND VGND VPWR VPWR _01941_ sky130_fd_sc_hd__or2_1
XFILLER_0_116_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_539 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07166_ net168 _01175_ VGND VGND VPWR VPWR _01186_ sky130_fd_sc_hd__and2b_1
XFILLER_0_112_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07097_ _00420_ VGND VGND VPWR VPWR _00431_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09273__A _01412_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09807_ _01995_ _01997_ VGND VGND VPWR VPWR _01998_ sky130_fd_sc_hd__or2_1
X_07999_ _02335_ _04917_ _04939_ _03070_ VGND VGND VPWR VPWR _00043_ sky130_fd_sc_hd__a22o_1
XANTENNA__12411__B _01584_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09738_ _00891_ _01545_ net52 _03587_ VGND VGND VPWR VPWR _01922_ sky130_fd_sc_hd__a22oi_1
XANTENNA__10212__A _00157_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09669_ _01844_ _01845_ VGND VGND VPWR VPWR _01846_ sky130_fd_sc_hd__nor2_1
XTAP_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11700_ _04068_ _04074_ VGND VGND VPWR VPWR _04075_ sky130_fd_sc_hd__xor2_1
XTAP_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12680_ _05141_ _05142_ _05144_ VGND VGND VPWR VPWR _05153_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_49_250 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11631_ _01155_ _01957_ _03951_ _03952_ VGND VGND VPWR VPWR _03999_ sky130_fd_sc_hd__a211o_1
XTAP_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12784__D _02849_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11562_ _03898_ _03903_ VGND VGND VPWR VPWR _03923_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10513_ _02768_ _02769_ VGND VGND VPWR VPWR _02770_ sky130_fd_sc_hd__nand2_1
X_13301_ _05743_ VGND VGND VPWR VPWR _05823_ sky130_fd_sc_hd__inv_2
X_11493_ _03811_ _03836_ _03837_ VGND VGND VPWR VPWR _03847_ sky130_fd_sc_hd__and3_1
XFILLER_0_135_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13232_ _02716_ _02713_ _02715_ _05579_ _05757_ VGND VGND VPWR VPWR _05758_ sky130_fd_sc_hd__a41o_1
X_10444_ _02424_ _02437_ VGND VGND VPWR VPWR _02695_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07894__C _06818_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13163_ _05465_ _03624_ _03490_ VGND VGND VPWR VPWR _05684_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_0_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10375_ _06819_ _00413_ _00571_ _06821_ VGND VGND VPWR VPWR _02619_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08071__B _00114_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12114_ _04522_ _04529_ VGND VGND VPWR VPWR _04530_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_103_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13094_ _03668_ _05607_ VGND VGND VPWR VPWR _05608_ sky130_fd_sc_hd__xnor2_2
X_12045_ _04452_ _04453_ VGND VGND VPWR VPWR _04454_ sky130_fd_sc_hd__xor2_4
XFILLER_0_46_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12602__A _00914_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09183__A _01312_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13996_ _06576_ _06568_ _06574_ VGND VGND VPWR VPWR _06583_ sky130_fd_sc_hd__nor3_1
XANTENNA__10479__D _02730_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12947_ _05446_ _04454_ VGND VGND VPWR VPWR _05447_ sky130_fd_sc_hd__xnor2_4
XANTENNA__09864__A1 _00004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13660__A2 _01958_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09864__B2 _07004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11671__A1 _07010_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11671__B2 _00101_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12878_ _01507_ _01369_ _01248_ _02117_ VGND VGND VPWR VPWR _05371_ sky130_fd_sc_hd__and4_1
XFILLER_0_56_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07431__A _04081_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11829_ _04165_ _02657_ _04166_ VGND VGND VPWR VPWR _04217_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_145_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07150__B _00989_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12620__B1 _01414_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12991__B _05483_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_130 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10792__A _05588_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09358__A _01368_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12215__C _00458_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08971_ _00969_ _01080_ VGND VGND VPWR VPWR _01082_ sky130_fd_sc_hd__and2_1
XFILLER_0_121_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07922_ _07045_ _07050_ VGND VGND VPWR VPWR _07051_ sky130_fd_sc_hd__xor2_1
X_07853_ net139 _06712_ _06939_ _06980_ VGND VGND VPWR VPWR _06982_ sky130_fd_sc_hd__o31ai_2
XANTENNA__09654__B1_N _01828_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07784_ _01044_ _00355_ _02960_ _03147_ VGND VGND VPWR VPWR _06913_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_824 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09523_ _01680_ _01685_ VGND VGND VPWR VPWR _01686_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09821__A _06819_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09454_ _01296_ _01294_ VGND VGND VPWR VPWR _01611_ sky130_fd_sc_hd__and2b_1
XFILLER_0_94_816 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07979__C _06819_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08405_ _00440_ _00462_ VGND VGND VPWR VPWR _00463_ sky130_fd_sc_hd__xnor2_1
X_09385_ _00459_ _01399_ _01534_ VGND VGND VPWR VPWR _01535_ sky130_fd_sc_hd__and3_1
XFILLER_0_59_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08336_ _03707_ VGND VGND VPWR VPWR _00389_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08267_ _00306_ _00307_ _00309_ _00312_ VGND VGND VPWR VPWR _00313_ sky130_fd_sc_hd__nor4_1
XFILLER_0_62_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_623 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07218_ _00442_ _00989_ _01744_ _00311_ VGND VGND VPWR VPWR _01755_ sky130_fd_sc_hd__and4_2
XFILLER_0_116_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08172__A _00208_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08198_ _00233_ _00241_ VGND VGND VPWR VPWR _00242_ sky130_fd_sc_hd__nand2_2
XFILLER_0_42_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07149_ net60 VGND VGND VPWR VPWR _01000_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_30_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10160_ _02382_ _02383_ VGND VGND VPWR VPWR _02384_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09715__B _00607_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10091_ _01350_ _02305_ _02307_ VGND VGND VPWR VPWR _02308_ sky130_fd_sc_hd__and3_2
XANTENNA__07516__A net6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11038__A net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13850_ _05907_ _05911_ _06421_ VGND VGND VPWR VPWR _06422_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_16_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12801_ _05106_ _05285_ VGND VGND VPWR VPWR _05286_ sky130_fd_sc_hd__nor2_1
X_10993_ _03270_ _03297_ VGND VGND VPWR VPWR _03298_ sky130_fd_sc_hd__nor2_1
X_13781_ _06334_ _06338_ _06345_ _06337_ VGND VGND VPWR VPWR _06346_ sky130_fd_sc_hd__o22a_1
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13253__A _05524_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12732_ _05169_ _05157_ _05158_ VGND VGND VPWR VPWR _05210_ sky130_fd_sc_hd__nand3_1
XANTENNA__08347__A _00344_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07251__A _02105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_743 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12663_ _05125_ _05128_ VGND VGND VPWR VPWR _05134_ sky130_fd_sc_hd__xor2_2
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11614_ _03974_ _03975_ _03976_ VGND VGND VPWR VPWR _03980_ sky130_fd_sc_hd__nand3_1
XFILLER_0_37_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09074__A2 _00423_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12594_ _05056_ _05057_ VGND VGND VPWR VPWR _05058_ sky130_fd_sc_hd__nor2_1
XFILLER_0_107_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11545_ _03898_ _03903_ VGND VGND VPWR VPWR _03904_ sky130_fd_sc_hd__or2b_1
XFILLER_0_108_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11476_ _03554_ _00508_ _01954_ _02135_ VGND VGND VPWR VPWR _03829_ sky130_fd_sc_hd__and4_1
XFILLER_0_123_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13215_ _05738_ _05739_ _05740_ VGND VGND VPWR VPWR _05741_ sky130_fd_sc_hd__a21oi_1
X_10427_ _02671_ _02676_ VGND VGND VPWR VPWR _02677_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14195_ _06636_ _06789_ VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__xor2_1
XANTENNA__10117__A _06937_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10358_ _07010_ _03685_ _00423_ _00101_ VGND VGND VPWR VPWR _02601_ sky130_fd_sc_hd__a22o_1
X_13146_ _05652_ _05653_ VGND VGND VPWR VPWR _05666_ sky130_fd_sc_hd__xnor2_1
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13077_ _02704_ _02705_ _02707_ VGND VGND VPWR VPWR _05590_ sky130_fd_sc_hd__a21oi_1
X_10289_ _05742_ _01545_ _02156_ _00628_ VGND VGND VPWR VPWR _02525_ sky130_fd_sc_hd__a22o_1
X_12028_ _04365_ _04435_ VGND VGND VPWR VPWR _04436_ sky130_fd_sc_hd__and2_1
XANTENNA__07426__A _04026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13979_ _05951_ _06156_ VGND VGND VPWR VPWR _06564_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07161__A _01120_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09170_ _01298_ _01299_ VGND VGND VPWR VPWR _01300_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08121_ _00156_ _00164_ VGND VGND VPWR VPWR _00165_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12507__A _04059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08704__B _00989_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08052_ _00497_ _00095_ VGND VGND VPWR VPWR _00096_ sky130_fd_sc_hd__nand2_1
XANTENNA__09088__A net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12226__B _01517_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09816__A _01188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08954_ _00775_ _00977_ _00976_ _00979_ VGND VGND VPWR VPWR _01063_ sky130_fd_sc_hd__o211a_1
XANTENNA__09535__B _02960_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07905_ _06970_ _07032_ _07006_ VGND VGND VPWR VPWR _07034_ sky130_fd_sc_hd__nand3_1
XANTENNA__10135__A1 _02971_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08885_ _00874_ _00876_ VGND VGND VPWR VPWR _00988_ sky130_fd_sc_hd__nor2_1
XANTENNA__10135__B2 _00366_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07836_ _06964_ VGND VGND VPWR VPWR _06965_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07767_ _06680_ _06701_ _06895_ VGND VGND VPWR VPWR _06896_ sky130_fd_sc_hd__nand3_1
X_09506_ _01665_ _01666_ VGND VGND VPWR VPWR _01668_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07698_ _06809_ _06816_ _06826_ VGND VGND VPWR VPWR _06827_ sky130_fd_sc_hd__and3_1
XFILLER_0_94_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09437_ _01583_ _01280_ _01590_ VGND VGND VPWR VPWR _01593_ sky130_fd_sc_hd__or3_1
XFILLER_0_109_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09368_ _00779_ VGND VGND VPWR VPWR _01517_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_47_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08319_ _00354_ _00368_ VGND VGND VPWR VPWR _00370_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09299_ _01440_ VGND VGND VPWR VPWR _01441_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11330_ _03654_ _03662_ VGND VGND VPWR VPWR _03669_ sky130_fd_sc_hd__xor2_2
XFILLER_0_22_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11261_ _03591_ _03592_ VGND VGND VPWR VPWR _03593_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13000_ _05496_ _05502_ _05504_ VGND VGND VPWR VPWR _05505_ sky130_fd_sc_hd__a21boi_2
XANTENNA__12363__A2 _00457_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10212_ _00157_ _02120_ _01966_ VGND VGND VPWR VPWR _02441_ sky130_fd_sc_hd__and3_1
X_11192_ _01156_ _01108_ _03515_ _03035_ VGND VGND VPWR VPWR _03517_ sky130_fd_sc_hd__a211o_1
X_10143_ _04862_ _00373_ _00782_ _04873_ VGND VGND VPWR VPWR _02365_ sky130_fd_sc_hd__a22oi_1
XANTENNA__14070__C _02743_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_394 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10074_ _02287_ _02288_ VGND VGND VPWR VPWR _02289_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13902_ _06453_ _06478_ VGND VGND VPWR VPWR _06479_ sky130_fd_sc_hd__and2_1
XANTENNA__12302__D _01505_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13833_ _06370_ _06381_ _06380_ VGND VGND VPWR VPWR _06403_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_134_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13764_ _06325_ _06326_ VGND VGND VPWR VPWR _06327_ sky130_fd_sc_hd__or2_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08077__A _06874_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10976_ _03258_ _03256_ VGND VGND VPWR VPWR _03280_ sky130_fd_sc_hd__and2b_1
XANTENNA__11215__B _03540_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12715_ _04691_ _05190_ VGND VGND VPWR VPWR _05191_ sky130_fd_sc_hd__nor2_2
XFILLER_0_85_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13695_ _02426_ _02737_ _06244_ VGND VGND VPWR VPWR _06251_ sky130_fd_sc_hd__and3_1
XFILLER_0_127_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12646_ _05108_ _05114_ VGND VGND VPWR VPWR _05116_ sky130_fd_sc_hd__xor2_1
XFILLER_0_143_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12577_ _00389_ _00393_ _01934_ _02169_ VGND VGND VPWR VPWR _05040_ sky130_fd_sc_hd__and4_1
XFILLER_0_108_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11528_ _03716_ _03885_ VGND VGND VPWR VPWR _03886_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10601__A2 _01410_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11459_ _03797_ _03809_ VGND VGND VPWR VPWR _03810_ sky130_fd_sc_hd__nor2_1
X_14178_ _06687_ _06777_ _06645_ VGND VGND VPWR VPWR _06778_ sky130_fd_sc_hd__a21oi_4
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13129_ _05644_ _05646_ VGND VGND VPWR VPWR _05647_ sky130_fd_sc_hd__xnor2_4
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07156__A _00869_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08670_ _05731_ net8 _03718_ _01000_ VGND VGND VPWR VPWR _00753_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09371__A _06483_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07621_ net140 _06120_ _06153_ VGND VGND VPWR VPWR _06164_ sky130_fd_sc_hd__a21o_1
XFILLER_0_108_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_440 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07552_ _03224_ _03235_ _03202_ VGND VGND VPWR VPWR _05423_ sky130_fd_sc_hd__o21ba_4
XANTENNA__11406__A _00257_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10310__A _00366_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07483_ _00661_ _04367_ VGND VGND VPWR VPWR _04664_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09222_ _01168_ _01165_ _01162_ VGND VGND VPWR VPWR _01357_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_146_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_746 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09153_ _01270_ _01217_ _01279_ VGND VGND VPWR VPWR _01281_ sky130_fd_sc_hd__and3_1
XFILLER_0_146_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_159 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08104_ _00045_ _00147_ VGND VGND VPWR VPWR _00148_ sky130_fd_sc_hd__nor2_1
XFILLER_0_126_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09084_ _00905_ _00908_ _01205_ VGND VGND VPWR VPWR _01206_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_140_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08035_ net165 _07075_ _00077_ VGND VGND VPWR VPWR _00079_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10980__A _00158_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11795__B _00159_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09986_ _02191_ _02192_ VGND VGND VPWR VPWR _02194_ sky130_fd_sc_hd__nor2_1
XANTENNA__07772__A2 _04851_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08937_ _00841_ _01043_ _01045_ VGND VGND VPWR VPWR _01046_ sky130_fd_sc_hd__o21a_2
X_08868_ _00797_ _00968_ VGND VGND VPWR VPWR _00970_ sky130_fd_sc_hd__or2_1
X_07819_ _06944_ _06947_ VGND VGND VPWR VPWR _06948_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09712__C _01508_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08799_ _00412_ _00562_ _00564_ VGND VGND VPWR VPWR _00895_ sky130_fd_sc_hd__nand3_1
XFILLER_0_39_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10830_ _04081_ net54 _02508_ _02507_ _02727_ VGND VGND VPWR VPWR _03119_ sky130_fd_sc_hd__a32o_1
XANTENNA__07513__B net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10220__A _05467_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07288__A1 _00891_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11035__B _01517_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10761_ _03011_ _03014_ _03006_ VGND VGND VPWR VPWR _03043_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_94_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12500_ _00612_ _03696_ _03729_ _04026_ VGND VGND VPWR VPWR _04955_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08047__D _06875_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13480_ _01108_ _03697_ _06011_ _06014_ VGND VGND VPWR VPWR _06015_ sky130_fd_sc_hd__o2bb2a_1
X_10692_ _00094_ _01411_ VGND VGND VPWR VPWR _02967_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12431_ _04777_ _04878_ VGND VGND VPWR VPWR _04879_ sky130_fd_sc_hd__nand2_1
XANTENNA__11689__C _00730_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12362_ _03696_ _03729_ net46 _01506_ VGND VGND VPWR VPWR _04803_ sky130_fd_sc_hd__and4_1
XFILLER_0_50_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10595__A1 _00310_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10595__B2 _00145_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14101_ _06612_ _06693_ _06694_ _05751_ VGND VGND VPWR VPWR _06696_ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07460__A1 _01470_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11313_ _03646_ _03648_ _03649_ VGND VGND VPWR VPWR _03650_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_132_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12293_ _00575_ _01664_ _01601_ _01505_ VGND VGND VPWR VPWR _04727_ sky130_fd_sc_hd__and4_1
XFILLER_0_31_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14032_ _06507_ _06607_ VGND VGND VPWR VPWR _06622_ sky130_fd_sc_hd__xnor2_4
X_11244_ _03569_ _03573_ VGND VGND VPWR VPWR _03574_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08360__A _00413_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11175_ _03470_ _03497_ VGND VGND VPWR VPWR _03498_ sky130_fd_sc_hd__xnor2_4
X_10126_ _02334_ _02345_ VGND VGND VPWR VPWR _02347_ sky130_fd_sc_hd__xnor2_1
X_10057_ _02151_ _02271_ VGND VGND VPWR VPWR _02272_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_54_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07704__A _01230_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13816_ _06374_ _06383_ VGND VGND VPWR VPWR _06385_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10130__A _00094_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13747_ _06300_ _06308_ VGND VGND VPWR VPWR _06309_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_512 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10959_ _00859_ _01400_ _03252_ _03251_ VGND VGND VPWR VPWR _03261_ sky130_fd_sc_hd__a31o_1
XFILLER_0_128_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13678_ _06074_ _06075_ _06177_ _06178_ VGND VGND VPWR VPWR _06233_ sky130_fd_sc_hd__a211o_1
XANTENNA__08535__A _00604_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13798__D _03680_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12629_ _05096_ _05086_ VGND VGND VPWR VPWR _05097_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_576 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13772__A1 _02765_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07203__A1 _00420_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10950__D _01504_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07203__B2 _00978_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09840_ _02031_ _02033_ VGND VGND VPWR VPWR _02034_ sky130_fd_sc_hd__xor2_1
XFILLER_0_95_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09771_ _01957_ VGND VGND VPWR VPWR _01958_ sky130_fd_sc_hd__buf_4
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08722_ _00808_ VGND VGND VPWR VPWR _00810_ sky130_fd_sc_hd__inv_2
X_08653_ net15 VGND VGND VPWR VPWR _00734_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__10510__A1 _01473_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07604_ _05654_ _05698_ _05665_ _05956_ VGND VGND VPWR VPWR _05977_ sky130_fd_sc_hd__a31o_1
XTAP_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08584_ _00653_ _00658_ VGND VGND VPWR VPWR _00659_ sky130_fd_sc_hd__and2b_1
XFILLER_0_76_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07535_ _04532_ _05225_ VGND VGND VPWR VPWR _05236_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_9_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10274__B1 net57 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12893__C _02133_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07466_ _04444_ _04466_ VGND VGND VPWR VPWR _04477_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_29_370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09205_ _01331_ _01336_ VGND VGND VPWR VPWR _01338_ sky130_fd_sc_hd__nor2_1
XFILLER_0_91_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07397_ net9 VGND VGND VPWR VPWR _03718_ sky130_fd_sc_hd__buf_4
XFILLER_0_134_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10026__B1 _01889_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09136_ _01194_ _01196_ _01259_ _01261_ VGND VGND VPWR VPWR _01263_ sky130_fd_sc_hd__o211a_1
XFILLER_0_72_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07442__A1 _03587_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09067_ _00416_ VGND VGND VPWR VPWR _01188_ sky130_fd_sc_hd__buf_4
XANTENNA__07442__B2 _03576_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08018_ _00059_ _00060_ net158 net171 VGND VGND VPWR VPWR _00062_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_102_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08942__A1 _00765_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09969_ _02167_ _02174_ VGND VGND VPWR VPWR _02175_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12980_ _04403_ _05482_ VGND VGND VPWR VPWR _05483_ sky130_fd_sc_hd__xor2_4
X_11931_ _00113_ _00114_ _00572_ _01272_ VGND VGND VPWR VPWR _04329_ sky130_fd_sc_hd__and4_1
XANTENNA__11691__D _01211_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11862_ _04142_ _04252_ VGND VGND VPWR VPWR _04253_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08058__C _00101_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13601_ _01414_ _03785_ _06136_ _06137_ VGND VGND VPWR VPWR _06148_ sky130_fd_sc_hd__o2bb2a_1
X_10813_ _03093_ _03098_ _03099_ VGND VGND VPWR VPWR _03100_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_67_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11793_ _04175_ _04176_ VGND VGND VPWR VPWR _04177_ sky130_fd_sc_hd__nor2_1
XFILLER_0_95_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13532_ _06059_ _06070_ VGND VGND VPWR VPWR _06072_ sky130_fd_sc_hd__or2_1
XFILLER_0_54_104 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10744_ _03017_ _03018_ _03020_ VGND VGND VPWR VPWR _03024_ sky130_fd_sc_hd__and3_1
XFILLER_0_94_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_796 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13463_ _01252_ _02737_ _05995_ VGND VGND VPWR VPWR _05996_ sky130_fd_sc_hd__a21boi_1
X_10675_ _02945_ _02947_ VGND VGND VPWR VPWR _02948_ sky130_fd_sc_hd__and2_1
XFILLER_0_125_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12414_ _04858_ _04859_ VGND VGND VPWR VPWR _04860_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13394_ _05915_ _05920_ VGND VGND VPWR VPWR _05921_ sky130_fd_sc_hd__and2_1
XFILLER_0_23_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_546 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12345_ _00915_ _01664_ VGND VGND VPWR VPWR _04784_ sky130_fd_sc_hd__nand2_1
XFILLER_0_121_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_732 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12276_ _04646_ _04702_ _04704_ VGND VGND VPWR VPWR _04709_ sky130_fd_sc_hd__nand3_1
XFILLER_0_121_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11866__D _00574_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14015_ _06599_ _06602_ VGND VGND VPWR VPWR _06603_ sky130_fd_sc_hd__xnor2_1
X_11227_ _03553_ _03555_ VGND VGND VPWR VPWR _03556_ sky130_fd_sc_hd__or2_1
XANTENNA__07418__B _03938_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output66_A net66 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11158_ _03478_ _03479_ VGND VGND VPWR VPWR _03480_ sky130_fd_sc_hd__xnor2_4
X_10109_ _02325_ _02327_ VGND VGND VPWR VPWR _02328_ sky130_fd_sc_hd__nor2_1
X_11089_ _03398_ _03403_ VGND VGND VPWR VPWR _03404_ sky130_fd_sc_hd__xnor2_4
XANTENNA__11882__C _02090_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12493__A1 _00374_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12245__A1 _00783_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10795__A _02259_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12245__B2 _04037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07320_ _02839_ _02861_ VGND VGND VPWR VPWR _02872_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08265__A _00298_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07251_ _02105_ VGND VGND VPWR VPWR _02116_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_73_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07182_ _01295_ VGND VGND VPWR VPWR _01361_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_54_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10019__B _04873_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12515__A _00374_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11776__D _01960_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10035__A _00859_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09823_ _06818_ _06820_ net9 net10 VGND VGND VPWR VPWR _02015_ sky130_fd_sc_hd__and4_1
X_09754_ _01917_ _01938_ VGND VGND VPWR VPWR _01939_ sky130_fd_sc_hd__xor2_2
X_08705_ _00431_ _04169_ net46 net47 VGND VGND VPWR VPWR _00791_ sky130_fd_sc_hd__and4_1
XANTENNA__12484__A1 _00374_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09685_ _01720_ _01485_ _01750_ _01749_ VGND VGND VPWR VPWR _01863_ sky130_fd_sc_hd__a31o_1
XFILLER_0_96_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10495__B1 _02731_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08636_ _00631_ _00715_ VGND VGND VPWR VPWR _00717_ sky130_fd_sc_hd__xnor2_1
XTAP_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08567_ _00637_ _00640_ VGND VGND VPWR VPWR _00641_ sky130_fd_sc_hd__and2_1
XFILLER_0_37_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07518_ _05016_ _05038_ VGND VGND VPWR VPWR _05049_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08498_ _00412_ _00564_ _00562_ VGND VGND VPWR VPWR _00566_ sky130_fd_sc_hd__a21oi_2
XANTENNA__07112__B1 net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12409__B _01584_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07449_ _04257_ _04279_ VGND VGND VPWR VPWR _04290_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_134_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10460_ _02711_ _02712_ VGND VGND VPWR VPWR _02713_ sky130_fd_sc_hd__nor2_4
XANTENNA__08903__A _00377_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09119_ _00344_ _01182_ _01229_ VGND VGND VPWR VPWR _01244_ sky130_fd_sc_hd__a21o_1
X_10391_ _02635_ _02636_ VGND VGND VPWR VPWR _02637_ sky130_fd_sc_hd__nand2_1
X_12130_ _04545_ _04547_ VGND VGND VPWR VPWR _04548_ sky130_fd_sc_hd__or2_4
XANTENNA__07966__A2 _07010_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12144__B _01183_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10970__A1 _04862_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10970__B2 _04873_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12061_ _04458_ _04465_ VGND VGND VPWR VPWR _04472_ sky130_fd_sc_hd__xor2_1
XFILLER_0_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09734__A _02467_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11012_ _03317_ _03318_ VGND VGND VPWR VPWR _03319_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12711__A2 _01062_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10722__A1 _01156_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07254__A _00650_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12963_ _04531_ _05463_ VGND VGND VPWR VPWR _05464_ sky130_fd_sc_hd__xor2_4
XANTENNA__09172__C _03707_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11914_ _04182_ _04206_ _04208_ _04309_ VGND VGND VPWR VPWR _04310_ sky130_fd_sc_hd__a211o_1
X_12894_ _05385_ _05386_ _05387_ VGND VGND VPWR VPWR _05388_ sky130_fd_sc_hd__a21oi_2
XANTENNA__07404__D _03718_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09891__A2 _02088_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12227__A1 _01517_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11845_ _04229_ _04233_ VGND VGND VPWR VPWR _04234_ sky130_fd_sc_hd__xor2_1
XFILLER_0_68_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output104_A net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12227__B2 _01518_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_142_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11776_ _05456_ _05478_ _02117_ _01960_ VGND VGND VPWR VPWR _04159_ sky130_fd_sc_hd__nand4_1
XTAP_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13515_ _06049_ _06052_ VGND VGND VPWR VPWR _06053_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_55_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10727_ _02994_ _03005_ VGND VGND VPWR VPWR _03006_ sky130_fd_sc_hd__xor2_1
XFILLER_0_83_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13446_ _05975_ _05976_ VGND VGND VPWR VPWR _05978_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10658_ _02769_ _02929_ VGND VGND VPWR VPWR _02930_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13377_ _01504_ _03738_ _03744_ _01508_ VGND VGND VPWR VPWR _05903_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10589_ _00310_ _01413_ _02844_ _02843_ VGND VGND VPWR VPWR _02854_ sky130_fd_sc_hd__a31o_1
XANTENNA__08532__B _02149_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10781__C _02725_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07957__A2 _00410_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07429__A _00442_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12328_ _01066_ _01188_ _03414_ _01289_ VGND VGND VPWR VPWR _04766_ sky130_fd_sc_hd__and4_1
XFILLER_0_23_398 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10961__A1 _00859_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08251__C _00293_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10961__B2 _01472_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12259_ _04688_ _04689_ VGND VGND VPWR VPWR _04690_ sky130_fd_sc_hd__xnor2_4
XANTENNA__10005__D _00613_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07590__B1 _00650_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12501__C _03685_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09470_ _01359_ _01425_ VGND VGND VPWR VPWR _01629_ sky130_fd_sc_hd__or2_1
XFILLER_0_92_89 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08421_ _00479_ _00480_ VGND VGND VPWR VPWR _00481_ sky130_fd_sc_hd__or2_1
XFILLER_0_116_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07893__A1 _00639_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07893__B2 net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10229__B1 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10956__C _01507_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08352_ _00401_ _00404_ _00405_ VGND VGND VPWR VPWR _00406_ sky130_fd_sc_hd__o21a_1
XFILLER_0_58_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12229__B _03750_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07303_ _00705_ net28 _00573_ net29 VGND VGND VPWR VPWR _02686_ sky130_fd_sc_hd__and4_1
XFILLER_0_129_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08283_ _00377_ _02982_ _06873_ _06874_ VGND VGND VPWR VPWR _00330_ sky130_fd_sc_hd__and4_1
XFILLER_0_144_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07234_ _01908_ _01919_ VGND VGND VPWR VPWR _01930_ sky130_fd_sc_hd__nand2_1
XFILLER_0_132_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07165_ _01022_ _01153_ VGND VGND VPWR VPWR _01175_ sky130_fd_sc_hd__nand2_1
XFILLER_0_131_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07096_ net1 VGND VGND VPWR VPWR _00420_ sky130_fd_sc_hd__buf_6
XFILLER_0_41_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09806_ _01981_ _01994_ VGND VGND VPWR VPWR _01997_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07998_ _07003_ _07036_ _00040_ VGND VGND VPWR VPWR _00042_ sky130_fd_sc_hd__a21oi_1
X_09737_ _04081_ _01410_ _01652_ _01651_ VGND VGND VPWR VPWR _01921_ sky130_fd_sc_hd__a31o_1
XFILLER_0_69_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10212__B _02120_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09668_ _00654_ _00859_ _01843_ VGND VGND VPWR VPWR _01845_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_139_404 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08619_ _00696_ _00697_ VGND VGND VPWR VPWR _00698_ sky130_fd_sc_hd__nor2_1
XFILLER_0_139_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09599_ _01765_ _01769_ VGND VGND VPWR VPWR _01770_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_84_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11630_ _03951_ _03952_ _01155_ _01958_ VGND VGND VPWR VPWR _03998_ sky130_fd_sc_hd__o211ai_1
XTAP_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_312 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11561_ _03919_ _03921_ VGND VGND VPWR VPWR _03922_ sky130_fd_sc_hd__and2b_1
XFILLER_0_119_172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13300_ _05713_ _05733_ VGND VGND VPWR VPWR _05822_ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10512_ _00636_ _01156_ _02765_ _02722_ VGND VGND VPWR VPWR _02769_ sky130_fd_sc_hd__and4_1
X_11492_ _03789_ _03845_ VGND VGND VPWR VPWR _03846_ sky130_fd_sc_hd__or2_1
XFILLER_0_33_630 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13231_ _05590_ _02711_ _05578_ VGND VGND VPWR VPWR _05757_ sky130_fd_sc_hd__o21a_1
XFILLER_0_134_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10443_ _02645_ _02693_ VGND VGND VPWR VPWR _02694_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_134_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07894__D net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13162_ _05669_ _05670_ VGND VGND VPWR VPWR _05683_ sky130_fd_sc_hd__xnor2_2
X_10374_ _06819_ _06821_ _00730_ VGND VGND VPWR VPWR _02618_ sky130_fd_sc_hd__and3_1
XFILLER_0_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12113_ _04523_ _04528_ VGND VGND VPWR VPWR _04529_ sky130_fd_sc_hd__xnor2_2
XANTENNA__14134__B2 _02743_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_595 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13093_ _03456_ _03496_ _03625_ _05606_ VGND VGND VPWR VPWR _05607_ sky130_fd_sc_hd__o31a_1
X_12044_ _04396_ _04397_ _04392_ VGND VGND VPWR VPWR _04453_ sky130_fd_sc_hd__o21bai_4
XANTENNA__12602__B _01412_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09561__A1 _00543_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09561__B2 _07040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09183__B _00543_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13995_ _05417_ _05954_ _05955_ _06580_ VGND VGND VPWR VPWR _06581_ sky130_fd_sc_hd__o211a_1
XFILLER_0_99_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13714__A _02426_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12946_ _05442_ _05443_ _05444_ VGND VGND VPWR VPWR _05446_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_62_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09864__A2 _00390_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08808__A _02127_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11671__A2 _00423_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12877_ _01507_ _02119_ VGND VGND VPWR VPWR _05370_ sky130_fd_sc_hd__nand2_1
XTAP_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11828_ _04150_ _04215_ VGND VGND VPWR VPWR _04216_ sky130_fd_sc_hd__xnor2_2
XANTENNA__07431__B _04048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07150__C _01000_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12620__A1 _01289_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11759_ _04124_ _04133_ VGND VGND VPWR VPWR _04140_ sky130_fd_sc_hd__nor2_1
XANTENNA__12620__B2 _01188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_602 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10792__B _01933_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13429_ _05851_ _05958_ _05959_ VGND VGND VPWR VPWR _05960_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_113_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08970_ _00969_ _01080_ VGND VGND VPWR VPWR _01081_ sky130_fd_sc_hd__nor2_1
X_07921_ _07048_ _07049_ VGND VGND VPWR VPWR _07050_ sky130_fd_sc_hd__nor2_1
X_07852_ net139 _06712_ _06939_ _06980_ VGND VGND VPWR VPWR _06981_ sky130_fd_sc_hd__or4_4
XANTENNA__10313__A _05203_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput1 a[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_4
X_07783_ _01044_ _03147_ _00355_ _02960_ VGND VGND VPWR VPWR _06912_ sky130_fd_sc_hd__and4_1
X_09522_ _01681_ _01684_ VGND VGND VPWR VPWR _01685_ sky130_fd_sc_hd__xor2_1
XFILLER_0_79_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09821__B _00423_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09453_ _01608_ _01609_ VGND VGND VPWR VPWR _01610_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_94_828 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07979__D _06821_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08404_ _00456_ _00461_ VGND VGND VPWR VPWR _00462_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_93_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09384_ _01532_ _01533_ VGND VGND VPWR VPWR _01534_ sky130_fd_sc_hd__xor2_1
XFILLER_0_47_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08335_ _00384_ _00386_ VGND VGND VPWR VPWR _00387_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08266_ _02280_ _00310_ _00308_ VGND VGND VPWR VPWR _00312_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_34_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_164 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07217_ _00672_ VGND VGND VPWR VPWR _01744_ sky130_fd_sc_hd__buf_4
XFILLER_0_132_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08197_ _00239_ _00240_ VGND VGND VPWR VPWR _00241_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07148_ _00978_ VGND VGND VPWR VPWR _00989_ sky130_fd_sc_hd__buf_4
XFILLER_0_70_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10090_ _01383_ _02306_ VGND VGND VPWR VPWR _02307_ sky130_fd_sc_hd__nand2_1
XANTENNA__11038__B _00373_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12800_ _05279_ _05284_ VGND VGND VPWR VPWR _05285_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13534__A _02766_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13780_ _06334_ _06344_ VGND VGND VPWR VPWR _06345_ sky130_fd_sc_hd__nor2_1
X_10992_ _03289_ _03295_ _03296_ VGND VGND VPWR VPWR _03297_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07532__A _05192_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12731_ _05157_ _05158_ _05169_ VGND VGND VPWR VPWR _05209_ sky130_fd_sc_hd__a21o_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08347__B _00391_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12662_ _04881_ _05036_ VGND VGND VPWR VPWR _05133_ sky130_fd_sc_hd__xor2_2
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11613_ _03829_ _03978_ VGND VGND VPWR VPWR _03979_ sky130_fd_sc_hd__nor2_1
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08806__B1 _00730_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12593_ _05054_ _05055_ _05053_ VGND VGND VPWR VPWR _05057_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_25_427 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09459__A net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11544_ _03901_ _03902_ VGND VGND VPWR VPWR _03903_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_80_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08363__A _00333_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11475_ _03814_ _03815_ VGND VGND VPWR VPWR _03827_ sky130_fd_sc_hd__xor2_1
X_13214_ _05682_ _05693_ VGND VGND VPWR VPWR _05740_ sky130_fd_sc_hd__and2_1
XFILLER_0_33_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10426_ _02672_ _02674_ VGND VGND VPWR VPWR _02676_ sky130_fd_sc_hd__xnor2_1
X_14194_ _06772_ _06773_ VGND VGND VPWR VPWR _06789_ sky130_fd_sc_hd__and2_1
XFILLER_0_21_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10117__B _02188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13145_ _05652_ _05653_ VGND VGND VPWR VPWR _05664_ sky130_fd_sc_hd__or2_1
X_10357_ _07010_ _00101_ _00423_ VGND VGND VPWR VPWR _02600_ sky130_fd_sc_hd__and3_1
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13076_ _05573_ VGND VGND VPWR VPWR _05589_ sky130_fd_sc_hd__inv_2
X_10288_ _00628_ _05742_ _01545_ VGND VGND VPWR VPWR _02524_ sky130_fd_sc_hd__and3_1
XANTENNA__09534__A1 _02971_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12027_ _04432_ _04434_ VGND VGND VPWR VPWR _04435_ sky130_fd_sc_hd__nor2_1
XANTENNA__09534__B2 _00366_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13978_ _05947_ _05952_ VGND VGND VPWR VPWR _06563_ sky130_fd_sc_hd__and2b_1
X_12929_ _04575_ _04580_ _04585_ VGND VGND VPWR VPWR _05427_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_76_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07161__B net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10852__B1 _02304_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08120_ _00162_ _00163_ VGND VGND VPWR VPWR _00164_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_83_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09369__A _00784_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12507__B _03938_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08704__C net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08051_ _00094_ VGND VGND VPWR VPWR _00095_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_114_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07784__B1 _02960_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08953_ _01061_ VGND VGND VPWR VPWR _01062_ sky130_fd_sc_hd__buf_4
X_07904_ _06970_ _07006_ _07032_ VGND VGND VPWR VPWR _07033_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_44_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08884_ _00874_ _00876_ VGND VGND VPWR VPWR _00987_ sky130_fd_sc_hd__nand2_1
XFILLER_0_138_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10135__A2 net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09832__A _07004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07835_ _06873_ VGND VGND VPWR VPWR _06964_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07766_ net150 _06175_ _06406_ _06615_ VGND VGND VPWR VPWR _06895_ sky130_fd_sc_hd__a211o_1
XFILLER_0_79_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09505_ _02116_ _02160_ _01508_ _01504_ VGND VGND VPWR VPWR _01666_ sky130_fd_sc_hd__and4_1
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07697_ _06824_ _06825_ VGND VGND VPWR VPWR _06826_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09436_ _01583_ _01280_ _01590_ VGND VGND VPWR VPWR _01592_ sky130_fd_sc_hd__o21ai_1
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09367_ _01382_ _01386_ VGND VGND VPWR VPWR _01516_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08318_ _00354_ _00368_ VGND VGND VPWR VPWR _00369_ sky130_fd_sc_hd__nor2_1
X_09298_ _01355_ _01163_ _01162_ VGND VGND VPWR VPWR _01440_ sky130_fd_sc_hd__or3b_2
XFILLER_0_35_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08249_ _00095_ VGND VGND VPWR VPWR _00293_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_105_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11260_ _03523_ _03527_ VGND VGND VPWR VPWR _03592_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_104_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10211_ _02115_ _02118_ _02121_ VGND VGND VPWR VPWR _02440_ sky130_fd_sc_hd__and3_1
X_11191_ _03515_ _03035_ _01156_ _01108_ VGND VGND VPWR VPWR _03516_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_101_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10142_ _02355_ _02363_ VGND VGND VPWR VPWR _02364_ sky130_fd_sc_hd__xnor2_2
XANTENNA__14070__D _02742_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10073_ _02256_ _02260_ _02286_ VGND VGND VPWR VPWR _02288_ sky130_fd_sc_hd__o21ai_1
X_13901_ _06465_ _06476_ _06477_ VGND VGND VPWR VPWR _06478_ sky130_fd_sc_hd__a21o_1
XANTENNA__13264__A _05507_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13832_ _06394_ _06399_ VGND VGND VPWR VPWR _06402_ sky130_fd_sc_hd__and2b_1
XANTENNA__09461__B _03894_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13763_ _06320_ _06322_ VGND VGND VPWR VPWR _06326_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10975_ _03276_ _03277_ VGND VGND VPWR VPWR _03278_ sky130_fd_sc_hd__nand2_1
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12714_ _00376_ _01183_ _01252_ _00380_ VGND VGND VPWR VPWR _05190_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_69_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13694_ _06243_ _06247_ _06249_ VGND VGND VPWR VPWR _06250_ sky130_fd_sc_hd__o21a_1
XFILLER_0_128_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12645_ _05111_ _05113_ VGND VGND VPWR VPWR _05114_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_127_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08805__B _04510_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09189__A _00257_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12576_ _04775_ net155 VGND VGND VPWR VPWR _05039_ sky130_fd_sc_hd__xor2_2
XFILLER_0_142_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_566 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11527_ _01312_ _01957_ _03690_ _01155_ VGND VGND VPWR VPWR _03885_ sky130_fd_sc_hd__a22oi_1
XANTENNA__11231__B _03559_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output96_A net96 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11458_ _03794_ _03796_ _03793_ VGND VGND VPWR VPWR _03809_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_111_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10409_ _02652_ _02656_ VGND VGND VPWR VPWR _02657_ sky130_fd_sc_hd__nand2_1
XANTENNA__13439__A _01181_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14177_ _05843_ _05849_ _06686_ VGND VGND VPWR VPWR _06777_ sky130_fd_sc_hd__a21o_1
X_11389_ _03723_ _03732_ VGND VGND VPWR VPWR _03733_ sky130_fd_sc_hd__and2b_1
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13128_ _05626_ _05645_ VGND VGND VPWR VPWR _05646_ sky130_fd_sc_hd__xnor2_4
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13303__A2 _05595_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13059_ _05565_ _05567_ _05569_ VGND VGND VPWR VPWR _05570_ sky130_fd_sc_hd__a21bo_1
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_46 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10798__A _06461_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07620_ _06098_ _06109_ VGND VGND VPWR VPWR _06153_ sky130_fd_sc_hd__and2_1
XANTENNA__09371__B _01517_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07551_ _05302_ _05401_ VGND VGND VPWR VPWR _05412_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11406__B _00670_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10310__B _02971_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10825__B1 net57 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07482_ _04400_ _04389_ VGND VGND VPWR VPWR _04653_ sky130_fd_sc_hd__or2b_1
XFILLER_0_146_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09221_ _01168_ _01169_ _01166_ VGND VGND VPWR VPWR _01356_ sky130_fd_sc_hd__and3_2
XFILLER_0_29_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_861 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07628__A2_N _05566_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_382 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09152_ _01270_ _01217_ _01279_ VGND VGND VPWR VPWR _01280_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_44_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_758 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08103_ _00141_ _00146_ VGND VGND VPWR VPWR _00147_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09083_ _00906_ _00907_ VGND VGND VPWR VPWR _01205_ sky130_fd_sc_hd__nand2_1
XFILLER_0_114_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10038__A _02246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08034_ _07039_ _07075_ _00077_ VGND VGND VPWR VPWR _00078_ sky130_fd_sc_hd__and3_1
XANTENNA__08731__A _00263_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10980__B _00457_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13349__A _01600_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11795__C _02459_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11553__A1 _06874_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07347__A _01044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11553__B2 _03510_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09985_ _06937_ _06637_ _02187_ _02189_ VGND VGND VPWR VPWR _02192_ sky130_fd_sc_hd__and4_1
XFILLER_0_110_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08936_ _00842_ _00872_ VGND VGND VPWR VPWR _01045_ sky130_fd_sc_hd__nand2_1
XANTENNA__07509__B1 _04939_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09562__A _00543_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08867_ _00797_ _00968_ VGND VGND VPWR VPWR _00969_ sky130_fd_sc_hd__nand2_1
X_07818_ _06945_ _06946_ VGND VGND VPWR VPWR _06947_ sky130_fd_sc_hd__xnor2_1
X_08798_ _00727_ _00893_ VGND VGND VPWR VPWR _00894_ sky130_fd_sc_hd__xnor2_2
XANTENNA__09712__D _01504_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07749_ _06824_ _06877_ VGND VGND VPWR VPWR _06878_ sky130_fd_sc_hd__xor2_2
XFILLER_0_67_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07513__C _04851_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10220__B _01000_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07288__A2 _01000_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10760_ _03031_ _03041_ VGND VGND VPWR VPWR _03042_ sky130_fd_sc_hd__and2b_1
XFILLER_0_67_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09419_ _01269_ _01282_ VGND VGND VPWR VPWR _01573_ sky130_fd_sc_hd__nand2_1
X_10691_ _02954_ _02953_ VGND VGND VPWR VPWR _02966_ sky130_fd_sc_hd__and2b_1
XANTENNA__08625__B _00703_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12430_ _04876_ _04877_ VGND VGND VPWR VPWR _04878_ sky130_fd_sc_hd__and2b_1
XFILLER_0_81_138 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11689__D net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12361_ _03729_ _00604_ _01506_ _03696_ VGND VGND VPWR VPWR _04802_ sky130_fd_sc_hd__a22o_1
XFILLER_0_117_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10595__A2 _02855_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14100_ _05648_ _05679_ _06694_ VGND VGND VPWR VPWR _06695_ sky130_fd_sc_hd__and3_1
X_11312_ _02913_ _03645_ VGND VGND VPWR VPWR _03649_ sky130_fd_sc_hd__nor2_1
XFILLER_0_133_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07460__A2 _04378_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12292_ _02187_ _01601_ _02189_ _00575_ VGND VGND VPWR VPWR _04726_ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14031_ _06598_ _06605_ VGND VGND VPWR VPWR _06621_ sky130_fd_sc_hd__xnor2_4
XANTENNA__09737__A1 _04081_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11243_ _03572_ _03560_ VGND VGND VPWR VPWR _03573_ sky130_fd_sc_hd__xor2_1
XFILLER_0_120_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11174_ _03471_ _03481_ VGND VGND VPWR VPWR _03497_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_101_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10125_ _02342_ _02344_ VGND VGND VPWR VPWR _02345_ sky130_fd_sc_hd__xnor2_2
X_10056_ _02242_ _02269_ VGND VGND VPWR VPWR _02271_ sky130_fd_sc_hd__xor2_2
XFILLER_0_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07704__B _00475_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13815_ _06366_ _06370_ _06372_ VGND VGND VPWR VPWR _06383_ sky130_fd_sc_hd__nor3_1
XANTENNA__10130__B _00784_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13746_ _06306_ _05872_ VGND VGND VPWR VPWR _06308_ sky130_fd_sc_hd__and2b_1
XFILLER_0_128_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10958_ _03255_ _03259_ VGND VGND VPWR VPWR _03260_ sky130_fd_sc_hd__or2b_1
XFILLER_0_57_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13677_ _06177_ _06178_ _06074_ _06075_ VGND VGND VPWR VPWR _06232_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_73_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10889_ _03182_ _03183_ VGND VGND VPWR VPWR _03184_ sky130_fd_sc_hd__nand2_1
X_12628_ _05094_ _05095_ VGND VGND VPWR VPWR _05096_ sky130_fd_sc_hd__xor2_1
XFILLER_0_109_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12559_ _05019_ _04975_ VGND VGND VPWR VPWR _05020_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_13_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14229_ _06810_ VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__inv_2
XFILLER_0_110_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07167__A net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07203__A2 _01208_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09770_ _01956_ VGND VGND VPWR VPWR _01957_ sky130_fd_sc_hd__clkbuf_4
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08721_ _00807_ _00808_ _00497_ _00142_ VGND VGND VPWR VPWR _00809_ sky130_fd_sc_hd__and4b_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08652_ _00731_ _00732_ VGND VGND VPWR VPWR _00733_ sky130_fd_sc_hd__or2b_1
XFILLER_0_96_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10510__A2 _02766_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07603_ _05709_ _05720_ _05956_ VGND VGND VPWR VPWR _05967_ sky130_fd_sc_hd__o21ai_2
X_08583_ _00655_ _00657_ VGND VGND VPWR VPWR _00658_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07534_ _01361_ _05181_ _05214_ VGND VGND VPWR VPWR _05225_ sky130_fd_sc_hd__and3_1
XFILLER_0_88_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10274__A1 _00989_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12893__D _02459_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10274__B2 _03576_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07465_ _00661_ _04455_ VGND VGND VPWR VPWR _04466_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12248__A _00379_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09204_ _01331_ _01336_ VGND VGND VPWR VPWR _01337_ sky130_fd_sc_hd__and2_1
XFILLER_0_91_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_579 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07396_ _03696_ VGND VGND VPWR VPWR _03707_ sky130_fd_sc_hd__buf_4
X_09135_ _05456_ _05478_ _03773_ _01260_ VGND VGND VPWR VPWR _01261_ sky130_fd_sc_hd__nand4_2
XANTENNA__07978__B1 _06821_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09557__A _00843_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09066_ _00940_ _00942_ _01185_ VGND VGND VPWR VPWR _01187_ sky130_fd_sc_hd__a21o_1
X_08017_ net159 _07061_ _00059_ _00060_ VGND VGND VPWR VPWR _00061_ sky130_fd_sc_hd__o211a_1
XFILLER_0_13_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13807__A _02190_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09968_ _02170_ _02173_ VGND VGND VPWR VPWR _02174_ sky130_fd_sc_hd__nand2_1
X_08919_ _00816_ _00834_ VGND VGND VPWR VPWR _01026_ sky130_fd_sc_hd__nand2_1
X_09899_ _02087_ _02097_ VGND VGND VPWR VPWR _02098_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11930_ _04324_ _04326_ _04327_ VGND VGND VPWR VPWR _04328_ sky130_fd_sc_hd__a21o_1
XANTENNA__10231__A _01306_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11861_ _04232_ _04251_ VGND VGND VPWR VPWR _04252_ sky130_fd_sc_hd__xnor2_2
X_13600_ _01061_ _03783_ _06146_ VGND VGND VPWR VPWR _06147_ sky130_fd_sc_hd__and3_1
XFILLER_0_39_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10812_ _03097_ _03095_ VGND VGND VPWR VPWR _03099_ sky130_fd_sc_hd__and2b_1
XFILLER_0_67_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08058__D _06733_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11792_ _02127_ net25 _04173_ _04174_ VGND VGND VPWR VPWR _04176_ sky130_fd_sc_hd__o2bb2a_1
X_13531_ _06059_ _06070_ VGND VGND VPWR VPWR _06071_ sky130_fd_sc_hd__nand2_1
XANTENNA__10265__A1 _00991_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10743_ _02886_ _03022_ VGND VGND VPWR VPWR _03023_ sky130_fd_sc_hd__or2_1
XANTENNA__11462__B1 _02133_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13462_ _05969_ _02735_ VGND VGND VPWR VPWR _05995_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10674_ _00294_ _02857_ _02946_ VGND VGND VPWR VPWR _02947_ sky130_fd_sc_hd__and3_1
XANTENNA__13203__A1 _05455_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12413_ _04841_ _04844_ VGND VGND VPWR VPWR _04859_ sky130_fd_sc_hd__xor2_1
X_13393_ _05916_ _05919_ VGND VGND VPWR VPWR _05920_ sky130_fd_sc_hd__xor2_1
XFILLER_0_106_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12344_ _04781_ _04778_ _04782_ VGND VGND VPWR VPWR _04783_ sky130_fd_sc_hd__and3_1
XFILLER_0_23_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_744 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12275_ _04637_ _04706_ VGND VGND VPWR VPWR _04707_ sky130_fd_sc_hd__nor2_1
X_14014_ _06502_ _06601_ VGND VGND VPWR VPWR _06602_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12714__B1 _01252_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11226_ _03234_ _03237_ _03232_ VGND VGND VPWR VPWR _03555_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_120_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07197__A1 _01284_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11157_ _03386_ _03402_ _03441_ _03384_ VGND VGND VPWR VPWR _03479_ sky130_fd_sc_hd__a31o_2
XANTENNA_max_cap130_A _05595_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10108_ _02323_ _01058_ _05577_ _02326_ VGND VGND VPWR VPWR _02327_ sky130_fd_sc_hd__and4b_1
X_11088_ _03396_ _03399_ VGND VGND VPWR VPWR _03403_ sky130_fd_sc_hd__nor2_2
XANTENNA__11882__D _01780_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10039_ _02250_ _02251_ VGND VGND VPWR VPWR _02252_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12493__A2 _00755_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12245__A2 _01178_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10795__B _02171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13729_ _06253_ _06288_ VGND VGND VPWR VPWR _06289_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07250_ _00628_ VGND VGND VPWR VPWR _02105_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_116_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07181_ _01339_ VGND VGND VPWR VPWR _01350_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_6_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10019__C _04037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12515__B _04059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10316__A _04598_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09822_ _06821_ net10 VGND VGND VPWR VPWR _02014_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07625__A _05467_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09753_ _01936_ _01937_ VGND VGND VPWR VPWR _01938_ sky130_fd_sc_hd__nand2_1
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08704_ _00442_ _00989_ net45 _00604_ VGND VGND VPWR VPWR _00790_ sky130_fd_sc_hd__and4_1
X_09684_ _01861_ VGND VGND VPWR VPWR _01862_ sky130_fd_sc_hd__inv_2
XFILLER_0_146_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12484__A2 _00741_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08635_ _00710_ _00714_ VGND VGND VPWR VPWR _00715_ sky130_fd_sc_hd__xnor2_2
XANTENNA__10495__A1 _00636_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10495__B2 _00526_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08566_ _00638_ VGND VGND VPWR VPWR _00640_ sky130_fd_sc_hd__inv_2
XTAP_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12236__A2 _03750_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07517_ _00300_ _05027_ VGND VGND VPWR VPWR _05038_ sky130_fd_sc_hd__nand2_1
XFILLER_0_147_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08497_ _00412_ _00562_ _00564_ VGND VGND VPWR VPWR _00565_ sky130_fd_sc_hd__and3_4
XFILLER_0_9_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07112__A1 _00563_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07112__B2 net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07448_ _04268_ _04048_ VGND VGND VPWR VPWR _04279_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07379_ _03510_ VGND VGND VPWR VPWR _03521_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_91_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08903__B _02993_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09118_ _01234_ _01237_ VGND VGND VPWR VPWR _01243_ sky130_fd_sc_hd__nor2b_4
XFILLER_0_44_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10390_ _02399_ _02409_ _02420_ VGND VGND VPWR VPWR _02636_ sky130_fd_sc_hd__o21ai_1
X_09049_ _01042_ _01046_ VGND VGND VPWR VPWR _01168_ sky130_fd_sc_hd__nand2_1
XFILLER_0_130_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10970__A2 _00604_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12060_ _04457_ _04470_ VGND VGND VPWR VPWR _04471_ sky130_fd_sc_hd__and2_1
X_11011_ _04598_ _00604_ VGND VGND VPWR VPWR _03318_ sky130_fd_sc_hd__nand2_1
XANTENNA__13537__A _03690_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09734__B _01060_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10722__A2 _02766_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13256__B _05779_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12962_ _05459_ _05461_ _05462_ VGND VGND VPWR VPWR _05463_ sky130_fd_sc_hd__or3_4
XANTENNA__09172__D _03740_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09750__A _00453_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11913_ _00157_ _00159_ _03683_ _03679_ VGND VGND VPWR VPWR _04309_ sky130_fd_sc_hd__and4_1
XFILLER_0_59_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12893_ _00783_ _00778_ _02133_ _02459_ VGND VGND VPWR VPWR _05387_ sky130_fd_sc_hd__and4_1
X_11844_ _04230_ _04227_ VGND VGND VPWR VPWR _04233_ sky130_fd_sc_hd__nand2_1
XTAP_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07270__A _00453_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11775_ _04151_ _04156_ VGND VGND VPWR VPWR _04157_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13514_ _06050_ _06051_ VGND VGND VPWR VPWR _06052_ sky130_fd_sc_hd__nand2_1
X_10726_ _02990_ _02991_ VGND VGND VPWR VPWR _03005_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13445_ _01183_ _01252_ _02766_ _02722_ VGND VGND VPWR VPWR _05976_ sky130_fd_sc_hd__and4_1
XFILLER_0_126_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10657_ _00636_ _02765_ _02722_ _01156_ VGND VGND VPWR VPWR _02929_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_125_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13376_ _00607_ _03744_ _05372_ _05371_ VGND VGND VPWR VPWR _05902_ sky130_fd_sc_hd__a31oi_2
X_10588_ _02847_ _02852_ VGND VGND VPWR VPWR _02853_ sky130_fd_sc_hd__or2b_1
XFILLER_0_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08532__C _04037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10781__D _02730_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12327_ _04762_ _04764_ VGND VGND VPWR VPWR _04765_ sky130_fd_sc_hd__xnor2_2
XANTENNA__07429__B _02051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10961__A2 _02188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08251__D _00294_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12258_ _00378_ _03738_ VGND VGND VPWR VPWR _04689_ sky130_fd_sc_hd__nand2_2
X_11209_ _03512_ _03534_ _03535_ VGND VGND VPWR VPWR _03536_ sky130_fd_sc_hd__o21a_1
XANTENNA__13447__A _01182_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12189_ _04611_ _04612_ VGND VGND VPWR VPWR _04613_ sky130_fd_sc_hd__or2_1
XANTENNA__07590__A1 _05456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07590__B2 _05467_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12501__D _00423_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_40 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08420_ _00478_ _00477_ VGND VGND VPWR VPWR _00480_ sky130_fd_sc_hd__and2b_1
XANTENNA__07893__A2 _06818_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07180__A _01230_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08351_ _00464_ _00381_ _00403_ VGND VGND VPWR VPWR _00405_ sky130_fd_sc_hd__a21o_1
XFILLER_0_19_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10956__D _01504_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10229__B2 _01470_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_723 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07302_ _02664_ _00672_ _00737_ _00726_ VGND VGND VPWR VPWR _02675_ sky130_fd_sc_hd__a31o_1
XFILLER_0_132_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08282_ _00254_ _00328_ VGND VGND VPWR VPWR _00329_ sky130_fd_sc_hd__xor2_1
XFILLER_0_132_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07233_ _01448_ _01832_ VGND VGND VPWR VPWR _01919_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_61_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07164_ _01022_ _01153_ VGND VGND VPWR VPWR _01164_ sky130_fd_sc_hd__nor2_1
XFILLER_0_131_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07095_ _00399_ VGND VGND VPWR VPWR _00410_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_140_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09090__A1_N _01744_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11692__A2_N _01211_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09805_ _01981_ _01994_ VGND VGND VPWR VPWR _01995_ sky130_fd_sc_hd__and2_1
X_07997_ _07003_ _07036_ _00040_ VGND VGND VPWR VPWR _00041_ sky130_fd_sc_hd__and3_1
X_09736_ _01654_ _01659_ VGND VGND VPWR VPWR _01920_ sky130_fd_sc_hd__nor2_1
X_09667_ _00654_ _00859_ _01843_ VGND VGND VPWR VPWR _01844_ sky130_fd_sc_hd__and3_1
XANTENNA__08530__B1 _02467_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08618_ _00505_ _00695_ VGND VGND VPWR VPWR _00697_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09598_ _01767_ _01768_ VGND VGND VPWR VPWR _01769_ sky130_fd_sc_hd__xnor2_1
XTAP_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07090__A net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08549_ _00619_ _00620_ VGND VGND VPWR VPWR _00621_ sky130_fd_sc_hd__or2_1
XTAP_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11560_ _03915_ _03920_ VGND VGND VPWR VPWR _03921_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10511_ _02764_ _02767_ VGND VGND VPWR VPWR _02768_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11491_ _03757_ _03782_ _03788_ VGND VGND VPWR VPWR _03845_ sky130_fd_sc_hd__and3_1
XFILLER_0_64_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11340__A _03678_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13230_ _02713_ _02714_ _05579_ VGND VGND VPWR VPWR _05756_ sky130_fd_sc_hd__and3_1
XFILLER_0_107_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10442_ _02690_ _02692_ VGND VGND VPWR VPWR _02693_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_123_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_686 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13161_ _05674_ _05681_ VGND VGND VPWR VPWR _05682_ sky130_fd_sc_hd__xor2_4
X_10373_ _02615_ _02616_ VGND VGND VPWR VPWR _02617_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12112_ _04525_ _04527_ VGND VGND VPWR VPWR _04528_ sky130_fd_sc_hd__xor2_4
XANTENNA__14134__A2 _02742_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13092_ _03672_ VGND VGND VPWR VPWR _05606_ sky130_fd_sc_hd__inv_2
X_12043_ _04406_ _04449_ _04450_ _04451_ VGND VGND VPWR VPWR _04452_ sky130_fd_sc_hd__o2bb2a_2
XANTENNA__07265__A _02259_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09561__A2 _01472_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09183__C _00636_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13994_ _06573_ _06579_ VGND VGND VPWR VPWR _06580_ sky130_fd_sc_hd__nor2_1
X_12945_ _04402_ _04471_ _04401_ VGND VGND VPWR VPWR _05444_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_87_314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13714__B _02759_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08521__B1 _00393_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08808__B _00734_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12876_ _01504_ _01249_ VGND VGND VPWR VPWR _05369_ sky130_fd_sc_hd__nand2_1
XTAP_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11827_ _04212_ _04214_ VGND VGND VPWR VPWR _04215_ sky130_fd_sc_hd__nor2_1
XTAP_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11959__A1 _06417_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11758_ _04126_ _04138_ VGND VGND VPWR VPWR _04139_ sky130_fd_sc_hd__xnor2_2
XANTENNA__07150__D _00901_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12620__A2 _01061_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10709_ _02959_ _02985_ VGND VGND VPWR VPWR _02986_ sky130_fd_sc_hd__or2_1
XFILLER_0_83_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_655 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_214 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12346__A _00916_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11689_ _06819_ _06821_ _00730_ net15 VGND VGND VPWR VPWR _04063_ sky130_fd_sc_hd__and4_1
XFILLER_0_3_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13428_ _05851_ _05957_ VGND VGND VPWR VPWR _05959_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13359_ _05867_ _05882_ VGND VGND VPWR VPWR _05883_ sky130_fd_sc_hd__xor2_1
XFILLER_0_140_157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07920_ _01000_ _04455_ _07046_ net173 VGND VGND VPWR VPWR _07049_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__07175__A _01076_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07851_ _06976_ _06979_ VGND VGND VPWR VPWR _06980_ sky130_fd_sc_hd__xor2_1
XANTENNA__10313__B _00604_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput2 a[10] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_2
X_07782_ _06909_ _06910_ VGND VGND VPWR VPWR _06911_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09521_ _01682_ _01683_ VGND VGND VPWR VPWR _01684_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_79_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09452_ _01285_ _01293_ _01286_ VGND VGND VPWR VPWR _01609_ sky130_fd_sc_hd__a21bo_1
X_08403_ _00453_ _00460_ VGND VGND VPWR VPWR _00461_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09383_ _06472_ _00458_ VGND VGND VPWR VPWR _01533_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08334_ _00385_ _00357_ VGND VGND VPWR VPWR _00386_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_52_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08265_ _00298_ VGND VGND VPWR VPWR _00310_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_46_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_817 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_491 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07216_ _01711_ _01722_ VGND VGND VPWR VPWR _01733_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08196_ _00234_ _00237_ _00236_ VGND VGND VPWR VPWR _00240_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_131_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07147_ net12 VGND VGND VPWR VPWR _00978_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_120_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07085__A net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10689__A1 _05203_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08909__A _06775_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09719_ _01672_ _01674_ _01899_ VGND VGND VPWR VPWR _01901_ sky130_fd_sc_hd__nor3_1
X_10991_ _03294_ _03292_ VGND VGND VPWR VPWR _03296_ sky130_fd_sc_hd__and2b_1
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12730_ _05196_ _05206_ _05207_ VGND VGND VPWR VPWR _05208_ sky130_fd_sc_hd__o21ai_4
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12661_ _04725_ _05131_ VGND VGND VPWR VPWR _05132_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_38_723 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11612_ _03554_ _01956_ _03687_ _00519_ VGND VGND VPWR VPWR _03978_ sky130_fd_sc_hd__a22oi_1
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12592_ _05053_ _05054_ _05055_ VGND VGND VPWR VPWR _05056_ sky130_fd_sc_hd__and3_1
XFILLER_0_53_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11543_ _03521_ _01960_ VGND VGND VPWR VPWR _03902_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09459__B _06820_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08363__B _00416_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11474_ _03823_ _03825_ VGND VGND VPWR VPWR _03826_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_122_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13213_ _05711_ _05696_ VGND VGND VPWR VPWR _05739_ sky130_fd_sc_hd__or2b_1
XFILLER_0_122_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10425_ _00322_ _02673_ VGND VGND VPWR VPWR _02674_ sky130_fd_sc_hd__nand2_1
XANTENNA__09231__A1 _01339_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14193_ _06641_ _06788_ VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14107__A2 _02742_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13144_ _05660_ _05662_ VGND VGND VPWR VPWR _05663_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_103_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10356_ _02397_ _02398_ VGND VGND VPWR VPWR _02599_ sky130_fd_sc_hd__and2_1
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13075_ _05563_ _05580_ _05586_ VGND VGND VPWR VPWR _05587_ sky130_fd_sc_hd__nand3_1
X_10287_ _02520_ _02522_ VGND VGND VPWR VPWR _02523_ sky130_fd_sc_hd__and2b_1
X_12026_ _04358_ _04362_ _04431_ VGND VGND VPWR VPWR _04434_ sky130_fd_sc_hd__nor3_1
XFILLER_0_73_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08819__A _00741_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07723__A _02105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13977_ _06547_ _06556_ _06561_ VGND VGND VPWR VPWR _06562_ sky130_fd_sc_hd__nor3_1
XFILLER_0_88_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12928_ _03613_ _05425_ VGND VGND VPWR VPWR _05426_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_76_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10852__A1 _03268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10852__B2 _05577_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12859_ _05273_ _05349_ VGND VGND VPWR VPWR _05350_ sky130_fd_sc_hd__or2_1
XFILLER_0_132_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10178__A2_N _03773_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08050_ _05203_ VGND VGND VPWR VPWR _00094_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_126_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08704__D _00604_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09385__A _00459_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07784__A1 _01044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08952_ _01060_ VGND VGND VPWR VPWR _01061_ sky130_fd_sc_hd__clkbuf_4
X_07903_ _07030_ _07031_ VGND VGND VPWR VPWR _07032_ sky130_fd_sc_hd__nor2_1
X_08883_ _00713_ _00985_ VGND VGND VPWR VPWR _00986_ sky130_fd_sc_hd__and2_1
XFILLER_0_37_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07834_ _06961_ _06962_ VGND VGND VPWR VPWR _06963_ sky130_fd_sc_hd__nor2_1
XANTENNA__09832__B _00390_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08729__A _00294_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07765_ _06883_ _06893_ VGND VGND VPWR VPWR _06894_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09504_ _02160_ _01664_ _01505_ _02116_ VGND VGND VPWR VPWR _01665_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_39_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07696_ _06822_ _06823_ _06817_ VGND VGND VPWR VPWR _06825_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_78_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09435_ _01588_ _01589_ VGND VGND VPWR VPWR _01590_ sky130_fd_sc_hd__and2_1
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10994__A _01473_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09366_ _01512_ _01513_ VGND VGND VPWR VPWR _01515_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__08464__A _00508_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08317_ net182 _00367_ VGND VGND VPWR VPWR _00368_ sky130_fd_sc_hd__xor2_2
X_09297_ _01431_ VGND VGND VPWR VPWR _01439_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08183__B _00219_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08248_ _00155_ _00154_ VGND VGND VPWR VPWR _00292_ sky130_fd_sc_hd__and2b_1
XFILLER_0_34_269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08179_ _00217_ _00219_ _00222_ VGND VGND VPWR VPWR _00223_ sky130_fd_sc_hd__a21o_1
XFILLER_0_132_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10210_ _02130_ _02140_ _02131_ VGND VGND VPWR VPWR _02439_ sky130_fd_sc_hd__a21bo_1
XANTENNA__07808__A _06472_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11190_ _03034_ VGND VGND VPWR VPWR _03515_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_820 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10141_ _02361_ _02362_ VGND VGND VPWR VPWR _02363_ sky130_fd_sc_hd__or2_2
X_10072_ _02256_ _02260_ _02286_ VGND VGND VPWR VPWR _02287_ sky130_fd_sc_hd__or3_1
X_13900_ _06463_ _06464_ _06457_ _06460_ VGND VGND VPWR VPWR _06477_ sky130_fd_sc_hd__o211a_1
X_13831_ _06392_ _06400_ VGND VGND VPWR VPWR _06401_ sky130_fd_sc_hd__nand2_1
XANTENNA__13264__B _05524_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09461__C _00475_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10974_ _04917_ _04939_ _00460_ _01400_ VGND VGND VPWR VPWR _03277_ sky130_fd_sc_hd__and4_1
X_13762_ _06277_ _06324_ VGND VGND VPWR VPWR _06325_ sky130_fd_sc_hd__and2_1
XFILLER_0_97_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12713_ _05184_ _05185_ _05188_ VGND VGND VPWR VPWR _05189_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_57_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14025__A1 _05810_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13693_ _06242_ _06248_ VGND VGND VPWR VPWR _06249_ sky130_fd_sc_hd__nor2_1
X_12644_ _05059_ _05083_ _05112_ VGND VGND VPWR VPWR _05113_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12587__A1 _00915_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08805__C net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09189__B _00670_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12575_ _04881_ _05036_ _04879_ VGND VGND VPWR VPWR _05037_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_92_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11526_ _03880_ _03882_ VGND VGND VPWR VPWR _03884_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11457_ _03801_ _03803_ _03807_ VGND VGND VPWR VPWR _03808_ sky130_fd_sc_hd__o21ai_2
XANTENNA__12624__A _00414_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10408_ _02654_ _02655_ VGND VGND VPWR VPWR _02656_ sky130_fd_sc_hd__xnor2_1
X_14176_ _06752_ _06759_ VGND VGND VPWR VPWR _06776_ sky130_fd_sc_hd__nor2_1
X_11388_ _03708_ _03731_ VGND VGND VPWR VPWR _03732_ sky130_fd_sc_hd__xor2_1
XANTENNA_output89_A net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13439__B _01250_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10339_ _02349_ _02375_ VGND VGND VPWR VPWR _02580_ sky130_fd_sc_hd__nand2_1
X_13127_ _05605_ _05623_ VGND VGND VPWR VPWR _05645_ sky130_fd_sc_hd__xnor2_2
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10144__A _04851_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13058_ _00381_ _00391_ VGND VGND VPWR VPWR _05569_ sky130_fd_sc_hd__nand2_2
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09933__A _02134_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12009_ _04413_ _04414_ VGND VGND VPWR VPWR _04415_ sky130_fd_sc_hd__nor2_1
XFILLER_0_84_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10798__B _02168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07550_ _05368_ _05390_ VGND VGND VPWR VPWR _05401_ sky130_fd_sc_hd__nor2_1
XANTENNA__07172__B net149 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11406__C _03750_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10310__C _01368_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10825__A1 _01339_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10825__B2 _04081_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07481_ _00300_ _04598_ _04631_ VGND VGND VPWR VPWR _04642_ sky130_fd_sc_hd__and3_1
XFILLER_0_76_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09220_ _01310_ _01353_ _01354_ VGND VGND VPWR VPWR _01355_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_119_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09151_ _01271_ _01278_ VGND VGND VPWR VPWR _01279_ sky130_fd_sc_hd__xor2_1
XFILLER_0_8_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09443__A1 _00416_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08102_ _02280_ _00145_ VGND VGND VPWR VPWR _00146_ sky130_fd_sc_hd__nand2_1
XFILLER_0_140_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09082_ _01202_ _01203_ VGND VGND VPWR VPWR _01204_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_364 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10038__B _02249_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08033_ _00075_ _00076_ VGND VGND VPWR VPWR _00077_ sky130_fd_sc_hd__xor2_2
XFILLER_0_114_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput60 b[5] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__buf_4
XFILLER_0_141_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08731__B _00819_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11002__A1 _05181_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13349__B _01585_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11795__D _02673_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11553__A2 _01177_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09984_ _06637_ _02188_ _02190_ _06937_ VGND VGND VPWR VPWR _02191_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_110_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08935_ _00842_ _00872_ VGND VGND VPWR VPWR _01043_ sky130_fd_sc_hd__nor2_1
XANTENNA__07509__A1 _00333_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08706__B1 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07509__B2 _02138_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12502__A1 _04048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09562__B _00859_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08866_ _00963_ _00966_ VGND VGND VPWR VPWR _00968_ sky130_fd_sc_hd__xor2_1
X_07817_ _02719_ net63 VGND VGND VPWR VPWR _06946_ sky130_fd_sc_hd__nand2_1
X_08797_ _00889_ _00892_ VGND VGND VPWR VPWR _00893_ sky130_fd_sc_hd__xnor2_2
X_07748_ _01350_ _06873_ _06876_ VGND VGND VPWR VPWR _06877_ sky130_fd_sc_hd__and3_1
XANTENNA__07513__D net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10220__C _01177_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07679_ _06755_ _06785_ VGND VGND VPWR VPWR _06790_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09418_ _01255_ _01571_ VGND VGND VPWR VPWR _01572_ sky130_fd_sc_hd__xnor2_4
X_10690_ _02961_ _02964_ VGND VGND VPWR VPWR _02965_ sky130_fd_sc_hd__or2b_1
XFILLER_0_75_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09349_ _05192_ net40 VGND VGND VPWR VPWR _01496_ sky130_fd_sc_hd__nand2_1
XANTENNA__09434__A1 _00157_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12360_ _04799_ _04800_ VGND VGND VPWR VPWR _04801_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_118_794 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11311_ _03635_ _03647_ VGND VGND VPWR VPWR _03648_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12291_ _04713_ _04724_ VGND VGND VPWR VPWR _04725_ sky130_fd_sc_hd__xor2_2
XFILLER_0_50_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14030_ _06619_ VGND VGND VPWR VPWR _06620_ sky130_fd_sc_hd__inv_2
XFILLER_0_132_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11242_ _03570_ _03571_ VGND VGND VPWR VPWR _03572_ sky130_fd_sc_hd__xnor2_2
XANTENNA__09737__A2 _01410_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11173_ _03490_ _03495_ VGND VGND VPWR VPWR _03496_ sky130_fd_sc_hd__and2_1
XFILLER_0_38_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10124_ _01912_ _01915_ _02203_ _02343_ VGND VGND VPWR VPWR _02344_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_100_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10055_ _02244_ _02268_ VGND VGND VPWR VPWR _02269_ sky130_fd_sc_hd__xnor2_4
XANTENNA_output127_A net127 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13814_ _06370_ _06380_ _06381_ VGND VGND VPWR VPWR _06382_ sky130_fd_sc_hd__or3_1
XFILLER_0_85_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13745_ _06301_ _06303_ _06305_ VGND VGND VPWR VPWR _06306_ sky130_fd_sc_hd__a21o_1
XFILLER_0_57_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10957_ _00145_ _00608_ _03256_ _03258_ VGND VGND VPWR VPWR _03259_ sky130_fd_sc_hd__a31o_1
XFILLER_0_97_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12619__A _00415_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07684__B1 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13676_ _06203_ _06229_ VGND VGND VPWR VPWR _06231_ sky130_fd_sc_hd__nor2_1
X_10888_ _03138_ _03167_ VGND VGND VPWR VPWR _03183_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11242__B _03571_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12627_ _01600_ _01060_ VGND VGND VPWR VPWR _05095_ sky130_fd_sc_hd__nand2_1
XANTENNA__10139__A _00457_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12558_ _04976_ _04967_ VGND VGND VPWR VPWR _05019_ sky130_fd_sc_hd__or2b_1
XFILLER_0_26_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11509_ _03863_ _03864_ VGND VGND VPWR VPWR _03865_ sky130_fd_sc_hd__and2_1
X_12489_ _01517_ _00916_ _04942_ VGND VGND VPWR VPWR _04943_ sky130_fd_sc_hd__and3_1
XFILLER_0_111_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07448__A _04268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14228_ _00244_ _00245_ _00242_ VGND VGND VPWR VPWR _06810_ sky130_fd_sc_hd__mux2_4
XFILLER_0_0_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14159_ _06698_ _06728_ VGND VGND VPWR VPWR _06759_ sky130_fd_sc_hd__or2_2
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_294 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09663__A _00670_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08720_ _03532_ _04895_ _04873_ _00121_ VGND VGND VPWR VPWR _00808_ sky130_fd_sc_hd__a22o_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07183__A _00891_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08651_ _01394_ net13 _00730_ _01470_ VGND VGND VPWR VPWR _00732_ sky130_fd_sc_hd__a22o_1
X_07602_ _05934_ _05945_ VGND VGND VPWR VPWR _05956_ sky130_fd_sc_hd__nor2_1
X_08582_ _00543_ _00656_ VGND VGND VPWR VPWR _00657_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07533_ _01405_ _05203_ VGND VGND VPWR VPWR _05214_ sky130_fd_sc_hd__nand2_1
XANTENNA__07911__A _04939_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09664__A1 _00843_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11471__A1 _00519_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07464_ net3 VGND VGND VPWR VPWR _04455_ sky130_fd_sc_hd__buf_2
XFILLER_0_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12248__B _03748_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09203_ _01332_ _01335_ VGND VGND VPWR VPWR _01336_ sky130_fd_sc_hd__xor2_1
XFILLER_0_119_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07395_ _03685_ VGND VGND VPWR VPWR _03696_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_146_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09134_ _03938_ VGND VGND VPWR VPWR _01260_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_45_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07978__A1 _00541_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07978__B2 net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09065_ _00740_ _00937_ _00936_ _00938_ VGND VGND VPWR VPWR _01185_ sky130_fd_sc_hd__o211a_1
XFILLER_0_130_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09557__B _00844_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08016_ _01197_ _04510_ net6 net7 VGND VGND VPWR VPWR _00060_ sky130_fd_sc_hd__nand4_1
XFILLER_0_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12723__A1 _00391_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09967_ _01934_ _02172_ VGND VGND VPWR VPWR _02173_ sky130_fd_sc_hd__nand2_1
X_08918_ _01007_ _01024_ VGND VGND VPWR VPWR _01025_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10512__A _00636_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09898_ _02095_ _02096_ VGND VGND VPWR VPWR _02097_ sky130_fd_sc_hd__nor2_1
XANTENNA__07093__A _00377_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08849_ _00947_ _00948_ VGND VGND VPWR VPWR _00949_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07524__C _00901_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10231__B _00672_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11860_ _04244_ _04247_ _04249_ _04250_ VGND VGND VPWR VPWR _04251_ sky130_fd_sc_hd__a31o_1
X_10811_ _03095_ _03097_ VGND VGND VPWR VPWR _03098_ sky130_fd_sc_hd__or2b_1
X_11791_ _04173_ _04174_ _01744_ net25 VGND VGND VPWR VPWR _04175_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_39_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09655__A1 _01626_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11343__A _03681_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13530_ _06068_ _06069_ VGND VGND VPWR VPWR _06070_ sky130_fd_sc_hd__nor2_1
XANTENNA__11462__A1 _00121_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10742_ _00635_ _01061_ _01414_ _07040_ VGND VGND VPWR VPWR _03022_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_94_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11462__B2 _03521_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10673_ _00293_ _02855_ VGND VGND VPWR VPWR _02946_ sky130_fd_sc_hd__nand2_1
X_13461_ _05969_ _02722_ _05980_ _05979_ VGND VGND VPWR VPWR _05994_ sky130_fd_sc_hd__a31o_1
XFILLER_0_137_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_448 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12412_ _04850_ _04856_ _04857_ VGND VGND VPWR VPWR _04858_ sky130_fd_sc_hd__a21o_1
XFILLER_0_35_353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09748__A net53 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13392_ _05917_ _05918_ VGND VGND VPWR VPWR _05919_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12343_ _01260_ _01506_ _01369_ _00755_ VGND VGND VPWR VPWR _04782_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12274_ _00376_ _01955_ _03686_ _00380_ VGND VGND VPWR VPWR _04706_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_10_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12714__A1 _00376_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14013_ _06501_ _06600_ VGND VGND VPWR VPWR _06601_ sky130_fd_sc_hd__nor2_1
X_11225_ _03232_ _03234_ _03237_ VGND VGND VPWR VPWR _03553_ sky130_fd_sc_hd__and3_1
XANTENNA__12714__B2 _00380_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07197__A2 _00672_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11156_ _03445_ _03476_ VGND VGND VPWR VPWR _03478_ sky130_fd_sc_hd__nand2_2
X_10107_ _05742_ net50 _01546_ _00628_ VGND VGND VPWR VPWR _02326_ sky130_fd_sc_hd__a22o_1
X_11087_ _03388_ _03396_ _03401_ VGND VGND VPWR VPWR _03402_ sky130_fd_sc_hd__or3_2
XANTENNA__08099__A _00142_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10038_ _02246_ _02249_ _01473_ _02247_ VGND VGND VPWR VPWR _02251_ sky130_fd_sc_hd__and4_1
XANTENNA__11237__B _03566_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07731__A _02664_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11989_ _03987_ VGND VGND VPWR VPWR _04393_ sky130_fd_sc_hd__inv_2
XANTENNA__12349__A _01260_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10795__C _02758_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13728_ _06250_ _06251_ VGND VGND VPWR VPWR _06288_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13659_ _06207_ _06209_ _06211_ VGND VGND VPWR VPWR _06212_ sky130_fd_sc_hd__a21o_1
XFILLER_0_38_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07180_ _01230_ VGND VGND VPWR VPWR _01339_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_90_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08562__A _04917_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10019__D _04059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08281__B _00327_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12515__C _03707_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10316__B net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09821_ _06819_ _00423_ VGND VGND VPWR VPWR _02013_ sky130_fd_sc_hd__nand2_1
X_09752_ _01932_ _01935_ VGND VGND VPWR VPWR _01937_ sky130_fd_sc_hd__or2_1
XANTENNA__07625__B _00541_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08703_ _00787_ _00788_ VGND VGND VPWR VPWR _00789_ sky130_fd_sc_hd__xnor2_2
X_09683_ _01859_ _01860_ VGND VGND VPWR VPWR _01861_ sky130_fd_sc_hd__nor2_1
XTAP_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08634_ _00251_ _00712_ _00713_ VGND VGND VPWR VPWR _00714_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10495__A2 _02735_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08565_ _03554_ _00508_ _04917_ _04939_ VGND VGND VPWR VPWR _00638_ sky130_fd_sc_hd__and4_1
XANTENNA__10247__A2 _02150_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07516_ net6 VGND VGND VPWR VPWR _05027_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_76_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11444__A1 _03554_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08496_ _04334_ _00348_ _04004_ VGND VGND VPWR VPWR _00564_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_119_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07112__A2 _00573_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07447_ _01230_ VGND VGND VPWR VPWR _04268_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_91_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07378_ _03499_ VGND VGND VPWR VPWR _03510_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_91_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09117_ _01239_ net131 VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__xnor2_4
XANTENNA__08903__C _00112_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10507__A _01472_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10955__B1 _01504_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09048_ _00877_ _00878_ _01047_ VGND VGND VPWR VPWR _01167_ sky130_fd_sc_hd__nor3_2
XANTENNA__07088__A _00322_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13818__A _01400_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12722__A _00380_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11010_ _03307_ _03306_ VGND VGND VPWR VPWR _03317_ sky130_fd_sc_hd__and2b_1
XFILLER_0_102_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09325__B1 _07040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12961_ _05444_ _05460_ VGND VGND VPWR VPWR _05462_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09750__B _01934_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11912_ _04161_ _04197_ _04199_ _04307_ VGND VGND VPWR VPWR _04308_ sky130_fd_sc_hd__a211o_1
XTAP_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12892_ _00784_ _02459_ VGND VGND VPWR VPWR _05386_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11843_ _04216_ _04231_ VGND VGND VPWR VPWR _04232_ sky130_fd_sc_hd__xnor2_2
XTAP_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07270__B _02280_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11774_ _04154_ _04155_ VGND VGND VPWR VPWR _04156_ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13513_ _05969_ _05985_ _02736_ _02737_ VGND VGND VPWR VPWR _06051_ sky130_fd_sc_hd__nand4_1
X_10725_ _03002_ VGND VGND VPWR VPWR _03003_ sky130_fd_sc_hd__inv_2
XTAP_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13444_ _05973_ _05974_ VGND VGND VPWR VPWR _05975_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10656_ _02924_ _02926_ VGND VGND VPWR VPWR _02928_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10587_ _00145_ _01413_ _02848_ _02851_ VGND VGND VPWR VPWR _02852_ sky130_fd_sc_hd__a31o_1
X_13375_ _05367_ _05374_ VGND VGND VPWR VPWR _05900_ sky130_fd_sc_hd__and2_1
XFILLER_0_51_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08532__D _04048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12326_ _00460_ _02090_ VGND VGND VPWR VPWR _04764_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07429__C _04037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12257_ _04676_ _04674_ VGND VGND VPWR VPWR _04688_ sky130_fd_sc_hd__or2b_2
XFILLER_0_76_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12632__A _00389_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output71_A net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11208_ _03498_ _03511_ VGND VGND VPWR VPWR _03535_ sky130_fd_sc_hd__or2_1
X_12188_ _03493_ _03622_ VGND VGND VPWR VPWR _04612_ sky130_fd_sc_hd__or2b_1
XANTENNA__13447__B _01252_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11139_ _03108_ _03248_ VGND VGND VPWR VPWR _03459_ sky130_fd_sc_hd__xor2_2
XANTENNA__07590__A2 _02105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09867__A1 _03521_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07461__A net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13182__B _05704_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08350_ _00464_ _00381_ _00403_ VGND VGND VPWR VPWR _00404_ sky130_fd_sc_hd__and3_1
XANTENNA__10229__A2 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07301_ net29 VGND VGND VPWR VPWR _02664_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_74_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08281_ _00290_ _00327_ VGND VGND VPWR VPWR _00328_ sky130_fd_sc_hd__xor2_2
XFILLER_0_58_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07232_ _01022_ _01897_ VGND VGND VPWR VPWR _01908_ sky130_fd_sc_hd__nand2_1
XANTENNA__11711__A _00257_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07163_ _01098_ _01142_ VGND VGND VPWR VPWR _01153_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_143_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07094_ _00388_ VGND VGND VPWR VPWR _00399_ sky130_fd_sc_hd__buf_4
XFILLER_0_14_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09804_ _01787_ _01993_ VGND VGND VPWR VPWR _01994_ sky130_fd_sc_hd__xnor2_1
X_07996_ _00038_ _00039_ VGND VGND VPWR VPWR _00040_ sky130_fd_sc_hd__xor2_1
X_09735_ _01339_ _01058_ _01657_ VGND VGND VPWR VPWR _01918_ sky130_fd_sc_hd__and3_1
XANTENNA__09570__B _01463_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09666_ _01840_ _01841_ VGND VGND VPWR VPWR _01843_ sky130_fd_sc_hd__nor2_1
XANTENNA__08467__A _02993_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08530__A1 _00453_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08530__B2 _00380_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08617_ _00505_ _00695_ VGND VGND VPWR VPWR _00696_ sky130_fd_sc_hd__and2_1
XTAP_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09597_ _00475_ net11 VGND VGND VPWR VPWR _01768_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08548_ _00444_ _00449_ _00618_ VGND VGND VPWR VPWR _00620_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_65_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08479_ _00399_ _00544_ VGND VGND VPWR VPWR _00545_ sky130_fd_sc_hd__nand2_1
XFILLER_0_108_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11621__A _00544_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10510_ _01473_ _02766_ _02761_ _02763_ VGND VGND VPWR VPWR _02767_ sky130_fd_sc_hd__a22oi_1
X_11490_ _03735_ _03843_ VGND VGND VPWR VPWR _03844_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10441_ _02142_ _02471_ _02691_ VGND VGND VPWR VPWR _02692_ sky130_fd_sc_hd__a21o_2
XFILLER_0_33_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09794__B1 _01600_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10372_ _02597_ _02395_ _02599_ _02614_ VGND VGND VPWR VPWR _02616_ sky130_fd_sc_hd__o31ai_2
X_13160_ _05668_ _05671_ VGND VGND VPWR VPWR _05681_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_33_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12111_ _04511_ _04513_ _04526_ VGND VGND VPWR VPWR _04527_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_32_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13091_ _04626_ _04627_ VGND VGND VPWR VPWR _05605_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_130_383 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12042_ _04407_ _04448_ VGND VGND VPWR VPWR _04451_ sky130_fd_sc_hd__nor2_1
XANTENNA__07265__B _00333_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09183__D _00526_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13993_ _05946_ _06563_ _06572_ VGND VGND VPWR VPWR _06579_ sky130_fd_sc_hd__nor3_1
X_12944_ _04581_ _04403_ VGND VGND VPWR VPWR _05443_ sky130_fd_sc_hd__nand2_1
XANTENNA__08521__A1 _03059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08521__B2 _02280_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12875_ _01180_ _05233_ _05235_ _05237_ VGND VGND VPWR VPWR _05367_ sky130_fd_sc_hd__o2bb2ai_1
XTAP_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11826_ _04193_ _04211_ VGND VGND VPWR VPWR _04214_ sky130_fd_sc_hd__and2_1
XTAP_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11959__A2 _02134_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11757_ _04132_ _04131_ VGND VGND VPWR VPWR _04138_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12627__A _01600_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10708_ _02956_ _02958_ VGND VGND VPWR VPWR _02985_ sky130_fd_sc_hd__nor2_1
XFILLER_0_83_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11688_ _03510_ _00734_ _02619_ _02618_ _00413_ VGND VGND VPWR VPWR _04062_ sky130_fd_sc_hd__a32o_1
XFILLER_0_126_667 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12346__B _01505_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13427_ _05417_ _05957_ VGND VGND VPWR VPWR _05958_ sky130_fd_sc_hd__xor2_2
X_10639_ _02862_ _02908_ VGND VGND VPWR VPWR _02909_ sky130_fd_sc_hd__xor2_1
XANTENNA__10919__B1 _02720_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13358_ _05880_ _05881_ VGND VGND VPWR VPWR _05882_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12309_ _04728_ _04732_ VGND VGND VPWR VPWR _04745_ sky130_fd_sc_hd__nor2_1
XANTENNA__12362__A _03696_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13289_ _05789_ _05807_ VGND VGND VPWR VPWR _05812_ sky130_fd_sc_hd__nand2_1
XFILLER_0_121_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07850_ _06883_ _06977_ _06978_ VGND VGND VPWR VPWR _06979_ sky130_fd_sc_hd__o21ai_1
X_07781_ _05060_ _06908_ VGND VGND VPWR VPWR _06910_ sky130_fd_sc_hd__and2_1
Xinput3 a[11] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_1
X_09520_ _01516_ _01520_ _01522_ _01385_ VGND VGND VPWR VPWR _01683_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_78_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09451_ _01596_ _01607_ VGND VGND VPWR VPWR _01608_ sky130_fd_sc_hd__xnor2_2
X_08402_ _00459_ VGND VGND VPWR VPWR _00460_ sky130_fd_sc_hd__buf_4
XFILLER_0_47_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09382_ _01530_ _01531_ VGND VGND VPWR VPWR _01532_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08333_ _00186_ _00249_ _00188_ _07083_ VGND VGND VPWR VPWR _00385_ sky130_fd_sc_hd__a31o_1
XFILLER_0_47_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08264_ _02040_ _00298_ _00308_ VGND VGND VPWR VPWR _00309_ sky130_fd_sc_hd__and3_1
XFILLER_0_116_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07215_ _01284_ _00300_ VGND VGND VPWR VPWR _01722_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08195_ _00238_ VGND VGND VPWR VPWR _00239_ sky130_fd_sc_hd__buf_2
XANTENNA__10057__A _02151_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07146_ _00912_ _00956_ VGND VGND VPWR VPWR _00967_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10504__B _07040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07979_ _00541_ _02719_ _06819_ _06821_ VGND VGND VPWR VPWR _00023_ sky130_fd_sc_hd__nand4_1
XANTENNA__08909__B _00151_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09718_ _01672_ _01674_ _01899_ VGND VGND VPWR VPWR _01900_ sky130_fd_sc_hd__o21a_1
XFILLER_0_69_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10990_ _03292_ _03294_ VGND VGND VPWR VPWR _03295_ sky130_fd_sc_hd__or2b_1
XFILLER_0_97_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09649_ _01822_ _01824_ VGND VGND VPWR VPWR _01825_ sky130_fd_sc_hd__xor2_4
XFILLER_0_97_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12660_ _05039_ _05130_ VGND VGND VPWR VPWR _05131_ sky130_fd_sc_hd__xnor2_1
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11611_ _03974_ _03975_ _03976_ VGND VGND VPWR VPWR _03977_ sky130_fd_sc_hd__a21o_1
XFILLER_0_38_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13260__B1 _05784_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12591_ _00745_ _02855_ _02857_ _00914_ VGND VGND VPWR VPWR _05055_ sky130_fd_sc_hd__a22o_1
XANTENNA__08806__A2 net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11542_ _03899_ _03900_ VGND VGND VPWR VPWR _03901_ sky130_fd_sc_hd__and2b_1
XFILLER_0_37_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09459__C net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11473_ _03808_ _03824_ VGND VGND VPWR VPWR _03825_ sky130_fd_sc_hd__and2_1
XFILLER_0_52_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13212_ _05682_ _05693_ VGND VGND VPWR VPWR _05738_ sky130_fd_sc_hd__or2_1
XFILLER_0_107_199 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09756__A _01889_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10424_ net25 VGND VGND VPWR VPWR _02673_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__08660__A _03773_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14192_ _06756_ _06757_ _06758_ VGND VGND VPWR VPWR _06788_ sky130_fd_sc_hd__and3_1
XFILLER_0_122_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09231__A2 _00604_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13143_ _05641_ _05661_ VGND VGND VPWR VPWR _05662_ sky130_fd_sc_hd__xnor2_4
X_10355_ _02065_ VGND VGND VPWR VPWR _02597_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10286_ _02159_ _02505_ _02506_ _02519_ VGND VGND VPWR VPWR _02522_ sky130_fd_sc_hd__a31o_1
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13074_ _02273_ _02491_ _02493_ _02713_ _05585_ VGND VGND VPWR VPWR _05586_ sky130_fd_sc_hd__a41o_1
XFILLER_0_57_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12025_ _04358_ _04362_ _04431_ VGND VGND VPWR VPWR _04432_ sky130_fd_sc_hd__o21a_1
XANTENNA__09491__A _00431_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07723__B _00650_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13976_ _06558_ _06559_ VGND VGND VPWR VPWR _06561_ sky130_fd_sc_hd__and2_1
X_12927_ _04617_ _04610_ VGND VGND VPWR VPWR _05425_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_860 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13741__A _02090_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10852__A2 _02158_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12858_ _05340_ _05348_ VGND VGND VPWR VPWR _05349_ sky130_fd_sc_hd__xor2_1
XTAP_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11809_ _04164_ _04170_ VGND VGND VPWR VPWR _04195_ sky130_fd_sc_hd__nor2_1
XTAP_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11899__C _03059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12789_ _05097_ _05272_ VGND VGND VPWR VPWR _05273_ sky130_fd_sc_hd__nor2_1
XTAP_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10605__A _00144_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07784__A2 _00355_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08951_ _01059_ VGND VGND VPWR VPWR _01060_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_121_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07902_ _07018_ _07029_ VGND VGND VPWR VPWR _07031_ sky130_fd_sc_hd__and2_1
X_08882_ _00710_ _00877_ VGND VGND VPWR VPWR _00985_ sky130_fd_sc_hd__nor2_1
XFILLER_0_138_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07914__A _00901_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07833_ _06870_ _06960_ VGND VGND VPWR VPWR _06962_ sky130_fd_sc_hd__and2_1
XANTENNA__11436__A _03750_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07764_ _06890_ _06892_ VGND VGND VPWR VPWR _06893_ sky130_fd_sc_hd__nor2_1
XANTENNA__09289__A2 _01233_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09503_ _01508_ VGND VGND VPWR VPWR _01664_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_78_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07695_ _06817_ _06822_ _06823_ VGND VGND VPWR VPWR _06824_ sky130_fd_sc_hd__and3_2
XFILLER_0_67_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09434_ _00157_ _01584_ _01587_ _01276_ VGND VGND VPWR VPWR _01589_ sky130_fd_sc_hd__a31o_1
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10994__B _02188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09365_ _01375_ _01378_ _01511_ VGND VGND VPWR VPWR _01513_ sky130_fd_sc_hd__nor3_1
XANTENNA__08464__B _00294_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08316_ _00358_ _00360_ _00362_ _00364_ _00365_ VGND VGND VPWR VPWR _00367_ sky130_fd_sc_hd__o311a_4
XFILLER_0_47_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09296_ _01433_ _01437_ VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__xor2_4
XFILLER_0_62_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08247_ _00156_ _00164_ VGND VGND VPWR VPWR _00291_ sky130_fd_sc_hd__nand2_1
XFILLER_0_117_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08178_ _00217_ _00219_ _00221_ VGND VGND VPWR VPWR _00222_ sky130_fd_sc_hd__o21ba_1
XANTENNA__10359__A1 _03696_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_432 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07129_ net29 net33 _00595_ _00584_ VGND VGND VPWR VPWR _00781_ sky130_fd_sc_hd__a31o_1
XFILLER_0_101_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__07096__A net1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10140_ _00458_ _02224_ _02360_ VGND VGND VPWR VPWR _02362_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_100_331 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10071_ _02284_ _02285_ VGND VGND VPWR VPWR _02286_ sky130_fd_sc_hd__nor2_1
XFILLER_0_100_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13545__B _02737_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13830_ _06394_ _06399_ VGND VGND VPWR VPWR _06400_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11346__A _02135_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13761_ _06268_ _06276_ VGND VGND VPWR VPWR _06324_ sky130_fd_sc_hd__or2_1
XANTENNA__12284__A1 _04714_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10973_ _03274_ _03275_ VGND VGND VPWR VPWR _03276_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12712_ _05183_ _05187_ VGND VGND VPWR VPWR _05188_ sky130_fd_sc_hd__nand2_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13692_ _02426_ _02736_ _02737_ _02427_ VGND VGND VPWR VPWR _06248_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_128_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12643_ _05052_ _05058_ VGND VGND VPWR VPWR _05112_ sky130_fd_sc_hd__and2b_1
XFILLER_0_38_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_811 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12587__A2 _01412_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08805__D _00730_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12574_ _04896_ _04910_ _05035_ _04893_ VGND VGND VPWR VPWR _05036_ sky130_fd_sc_hd__a31o_1
XFILLER_0_108_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09189__C _00819_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11525_ _03865_ _03881_ VGND VGND VPWR VPWR _03882_ sky130_fd_sc_hd__or2_1
XFILLER_0_80_343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11456_ _03804_ _03805_ VGND VGND VPWR VPWR _03807_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_80_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12624__B _00572_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10407_ _02029_ _01960_ VGND VGND VPWR VPWR _02655_ sky130_fd_sc_hd__nand2_1
X_14175_ _06771_ _06774_ VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__xnor2_1
XANTENNA__08412__B1 _00268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11387_ _03728_ _03730_ VGND VGND VPWR VPWR _03731_ sky130_fd_sc_hd__nor2_1
XFILLER_0_68_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10425__A _00322_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13439__C _02721_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13126_ _05639_ _05641_ _05642_ VGND VGND VPWR VPWR _05644_ sky130_fd_sc_hd__a21o_2
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10338_ _02545_ _02578_ VGND VGND VPWR VPWR _02579_ sky130_fd_sc_hd__xor2_4
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10144__B net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13057_ _05565_ _05567_ VGND VGND VPWR VPWR _05568_ sky130_fd_sc_hd__or2_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10269_ _02311_ _02320_ _02331_ VGND VGND VPWR VPWR _02503_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_84_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12640__A _00915_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12008_ _04329_ _04333_ _04412_ VGND VGND VPWR VPWR _04414_ sky130_fd_sc_hd__nor3_1
XANTENNA__09912__B1 _01249_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13959_ _06524_ _06525_ VGND VGND VPWR VPWR _06542_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11406__D _03748_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07480_ net33 _04367_ _04609_ _04620_ VGND VGND VPWR VPWR _04631_ sky130_fd_sc_hd__a31o_1
XANTENNA__08565__A _03554_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09150_ _01276_ _01277_ VGND VGND VPWR VPWR _01278_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10589__A1 _00310_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08101_ _00144_ VGND VGND VPWR VPWR _00145_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_71_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09081_ _00929_ _01201_ VGND VGND VPWR VPWR _01203_ sky130_fd_sc_hd__or2_1
XANTENNA__08651__B1 _00730_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10038__C _01473_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08032_ _07041_ _07073_ _07072_ VGND VGND VPWR VPWR _00076_ sky130_fd_sc_hd__a21o_1
XFILLER_0_71_376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput50 b[25] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_25_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput61 b[6] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_12_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11002__A2 _00604_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13349__C _02306_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07347__C _00880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09983_ _02189_ VGND VGND VPWR VPWR _02190_ sky130_fd_sc_hd__clkbuf_4
X_08934_ _01032_ _01041_ VGND VGND VPWR VPWR _01042_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_110_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08706__A1 _03587_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07509__A2 _04917_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08706__B2 _00431_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07644__A _05456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12502__A2 _03894_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08865_ _00964_ _00965_ VGND VGND VPWR VPWR _00966_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08182__A2 _03609_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07816_ net29 net63 _06858_ _06857_ VGND VGND VPWR VPWR _06945_ sky130_fd_sc_hd__a31o_1
X_08796_ _00631_ _00715_ _00890_ VGND VGND VPWR VPWR _00892_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_98_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07747_ _01383_ _06875_ VGND VGND VPWR VPWR _06876_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07678_ _00442_ _06765_ _06775_ _02051_ VGND VGND VPWR VPWR _06785_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_66_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14196__B _06778_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09417_ _01568_ _01570_ VGND VGND VPWR VPWR _01571_ sky130_fd_sc_hd__or2_2
XANTENNA__08890__B1 _04928_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09348_ _00612_ _01363_ _01494_ VGND VGND VPWR VPWR _01495_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_35_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09434__A2 _01584_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11777__B1 _01960_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09279_ _01417_ _01419_ VGND VGND VPWR VPWR _01420_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_708 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11310_ _02770_ _02787_ VGND VGND VPWR VPWR _03647_ sky130_fd_sc_hd__and2_1
XFILLER_0_90_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12290_ _04721_ _04723_ VGND VGND VPWR VPWR _04724_ sky130_fd_sc_hd__nor2_1
XFILLER_0_132_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11241_ _03419_ _03438_ VGND VGND VPWR VPWR _03571_ sky130_fd_sc_hd__xor2_4
X_11172_ _03494_ VGND VGND VPWR VPWR _03495_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10123_ _01904_ _01910_ _02202_ VGND VGND VPWR VPWR _02343_ sky130_fd_sc_hd__o21a_1
XFILLER_0_100_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10054_ _02266_ _02267_ VGND VGND VPWR VPWR _02268_ sky130_fd_sc_hd__nand2_2
XANTENNA__07554__A _01044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13813_ _03414_ _03679_ _06369_ VGND VGND VPWR VPWR _06381_ sky130_fd_sc_hd__a21oi_1
X_13744_ _05875_ _05881_ _06304_ VGND VGND VPWR VPWR _06305_ sky130_fd_sc_hd__o21a_1
XFILLER_0_58_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10956_ _04895_ _04873_ _01507_ _01504_ VGND VGND VPWR VPWR _03258_ sky130_fd_sc_hd__and4_1
XFILLER_0_97_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12619__B _00575_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07684__A1 net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13675_ _06220_ _06226_ _06228_ _06217_ VGND VGND VPWR VPWR _06229_ sky130_fd_sc_hd__o31a_1
XANTENNA__07684__B2 net149 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10887_ _03178_ _03181_ VGND VGND VPWR VPWR _03182_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12626_ _01413_ _05091_ _05092_ VGND VGND VPWR VPWR _05094_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_66_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12557_ _05014_ _05017_ VGND VGND VPWR VPWR _05018_ sky130_fd_sc_hd__xor2_4
XFILLER_0_79_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12635__A _00915_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11508_ _03835_ _03834_ VGND VGND VPWR VPWR _03864_ sky130_fd_sc_hd__xnor2_1
X_12488_ _01518_ _00914_ VGND VGND VPWR VPWR _04942_ sky130_fd_sc_hd__nand2_1
X_14227_ _00233_ _00241_ VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__xor2_1
X_11439_ _03754_ _03787_ VGND VGND VPWR VPWR _03788_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07448__B _04048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14158_ _05965_ _06754_ VGND VGND VPWR VPWR _06758_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13109_ _05217_ _05216_ VGND VGND VPWR VPWR _05625_ sky130_fd_sc_hd__or2b_1
XFILLER_0_0_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09663__B _00145_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14089_ _06649_ _06683_ VGND VGND VPWR VPWR _06684_ sky130_fd_sc_hd__xnor2_4
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08650_ _04510_ _00661_ net13 _00730_ VGND VGND VPWR VPWR _00731_ sky130_fd_sc_hd__and4_1
X_07601_ _05808_ _05923_ VGND VGND VPWR VPWR _05945_ sky130_fd_sc_hd__and2_1
X_08581_ _00388_ _02993_ _06765_ VGND VGND VPWR VPWR _00656_ sky130_fd_sc_hd__and3_1
XFILLER_0_88_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07532_ _05192_ VGND VGND VPWR VPWR _05203_ sky130_fd_sc_hd__buf_4
XFILLER_0_146_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07463_ _04422_ _04433_ VGND VGND VPWR VPWR _04444_ sky130_fd_sc_hd__and2b_1
XANTENNA__11471__A2 _03679_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09202_ _01333_ _01334_ VGND VGND VPWR VPWR _01335_ sky130_fd_sc_hd__or2_1
XFILLER_0_146_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07394_ net8 VGND VGND VPWR VPWR _03685_ sky130_fd_sc_hd__buf_6
XFILLER_0_91_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09133_ _05456_ _03773_ _03938_ _05467_ VGND VGND VPWR VPWR _01259_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07978__A2 _06818_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09064_ _00344_ _01183_ VGND VGND VPWR VPWR _01184_ sky130_fd_sc_hd__nand2_2
XFILLER_0_114_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08015_ _01197_ net6 net7 _01208_ VGND VGND VPWR VPWR _00059_ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_798 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12723__A2 _01062_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07920__A1_N _01000_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09966_ _03576_ _00989_ net54 VGND VGND VPWR VPWR _02172_ sky130_fd_sc_hd__and3_1
XFILLER_0_110_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08917_ _01020_ _01023_ VGND VGND VPWR VPWR _01024_ sky130_fd_sc_hd__xor2_1
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09897_ _02089_ _02093_ VGND VGND VPWR VPWR _02096_ sky130_fd_sc_hd__nor2_1
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10512__B _01156_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08848_ _05577_ _04026_ VGND VGND VPWR VPWR _00948_ sky130_fd_sc_hd__nand2_1
XANTENNA__07524__D _04378_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10231__C net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08779_ _00842_ _00872_ VGND VGND VPWR VPWR _00873_ sky130_fd_sc_hd__xnor2_1
X_10810_ _03063_ _03096_ VGND VGND VPWR VPWR _03097_ sky130_fd_sc_hd__nand2_1
X_11790_ _01295_ _02133_ net24 _01306_ VGND VGND VPWR VPWR _04174_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_138_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10741_ _03017_ _03018_ _03020_ VGND VGND VPWR VPWR _03021_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11462__A2 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_800 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13460_ _05986_ _05984_ VGND VGND VPWR VPWR _05993_ sky130_fd_sc_hd__or2b_1
XFILLER_0_48_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10672_ _02942_ _02943_ _02944_ VGND VGND VPWR VPWR _02945_ sky130_fd_sc_hd__and3_1
XFILLER_0_47_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12411_ _00378_ _01584_ _04854_ VGND VGND VPWR VPWR _04857_ sky130_fd_sc_hd__and3_1
XFILLER_0_36_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13391_ _01518_ _01517_ _03681_ _02673_ VGND VGND VPWR VPWR _05918_ sky130_fd_sc_hd__nand4_1
XFILLER_0_51_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12342_ _01260_ _00605_ _04779_ _04780_ VGND VGND VPWR VPWR _04781_ sky130_fd_sc_hd__a31o_1
XFILLER_0_105_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12273_ _04646_ _04702_ _04704_ VGND VGND VPWR VPWR _04705_ sky130_fd_sc_hd__a21o_1
X_14012_ _06499_ _06500_ VGND VGND VPWR VPWR _06600_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11224_ _03548_ _03549_ _02382_ _02588_ VGND VGND VPWR VPWR _03552_ sky130_fd_sc_hd__a211o_1
XANTENNA__09304__A_N _01311_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12714__A2 _01183_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11155_ _03443_ _03369_ VGND VGND VPWR VPWR _03476_ sky130_fd_sc_hd__nand2_1
XANTENNA__10703__A _00388_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07284__A _02456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10106_ _05588_ _01058_ _02322_ _02323_ VGND VGND VPWR VPWR _02325_ sky130_fd_sc_hd__o2bb2a_1
X_11086_ _03398_ _03399_ VGND VGND VPWR VPWR _03401_ sky130_fd_sc_hd__nor2_1
X_10037_ _02246_ _01473_ _02247_ _02249_ VGND VGND VPWR VPWR _02250_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_81_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07731__B _00475_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_12 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11988_ _04388_ _04390_ _04391_ VGND VGND VPWR VPWR _04392_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12349__B _00605_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10795__D _02169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13727_ _06284_ _06286_ VGND VGND VPWR VPWR _06287_ sky130_fd_sc_hd__and2b_1
X_10939_ _03232_ _03234_ _03237_ _03238_ VGND VGND VPWR VPWR _03239_ sky130_fd_sc_hd__a31o_1
XFILLER_0_58_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13658_ _06166_ _06210_ VGND VGND VPWR VPWR _06211_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_332 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12609_ _00915_ _01059_ VGND VGND VPWR VPWR _05075_ sky130_fd_sc_hd__nand2_1
XFILLER_0_144_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13589_ _06125_ _06134_ VGND VGND VPWR VPWR _06135_ sky130_fd_sc_hd__or2_1
XFILLER_0_5_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_516 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07459__A net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12953__A2 _05451_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12515__D _03740_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09820_ _03696_ _01761_ _01763_ _01764_ VGND VGND VPWR VPWR _02012_ sky130_fd_sc_hd__o2bb2ai_1
X_09751_ _01932_ _01935_ VGND VGND VPWR VPWR _01936_ sky130_fd_sc_hd__nand2_1
X_08702_ _00621_ _00622_ _00619_ VGND VGND VPWR VPWR _00788_ sky130_fd_sc_hd__o21bai_2
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09682_ _01857_ _01858_ VGND VGND VPWR VPWR _01860_ sky130_fd_sc_hd__nor2_1
XFILLER_0_146_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08633_ _00555_ _00711_ _00551_ VGND VGND VPWR VPWR _00713_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_12_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08564_ _00519_ _00636_ _00526_ _03554_ VGND VGND VPWR VPWR _00637_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07515_ _04994_ _05005_ VGND VGND VPWR VPWR _05016_ sky130_fd_sc_hd__or2b_1
X_08495_ _00439_ _00561_ VGND VGND VPWR VPWR _00562_ sky130_fd_sc_hd__xnor2_2
XANTENNA__11444__A2 _03678_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_654 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07446_ _01284_ net40 _04125_ _04114_ VGND VGND VPWR VPWR _04257_ sky130_fd_sc_hd__a31o_1
XFILLER_0_146_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__08753__A _00670_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07377_ net64 VGND VGND VPWR VPWR _03499_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_146_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09116_ _00894_ _00896_ _01054_ _01240_ _01053_ VGND VGND VPWR VPWR _01242_ sky130_fd_sc_hd__o32ai_2
XFILLER_0_44_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08903__D _00268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10955__A1 _04895_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10507__B _02759_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10955__B2 _04928_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09047_ _01162_ _01165_ VGND VGND VPWR VPWR _01166_ sky130_fd_sc_hd__and2_1
XFILLER_0_142_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09584__A _01486_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13818__B _02187_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12722__B _01182_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09949_ _01917_ _01936_ _01937_ VGND VGND VPWR VPWR _02153_ sky130_fd_sc_hd__a21bo_1
XANTENNA__09325__A1 _00654_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09325__B2 _00844_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12960_ _05436_ _05439_ _05441_ _05443_ _05460_ VGND VGND VPWR VPWR _05461_ sky130_fd_sc_hd__a311oi_4
X_11911_ _06626_ _06450_ _03750_ _03783_ VGND VGND VPWR VPWR _04307_ sky130_fd_sc_hd__and4_1
XTAP_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12891_ _00779_ _02134_ VGND VGND VPWR VPWR _05385_ sky130_fd_sc_hd__nand2_1
XTAP_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11842_ _04227_ _04229_ _04230_ VGND VGND VPWR VPWR _04231_ sky130_fd_sc_hd__a21bo_1
XTAP_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11773_ _01996_ _01960_ _04152_ _04153_ VGND VGND VPWR VPWR _04155_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_138_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13512_ _05985_ _02736_ _02737_ _05969_ VGND VGND VPWR VPWR _06050_ sky130_fd_sc_hd__a22o_1
XTAP_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10724_ _02935_ _03001_ VGND VGND VPWR VPWR _03002_ sky130_fd_sc_hd__xor2_1
XFILLER_0_83_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08663__A _00741_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13443_ _05969_ _02766_ _05971_ _05972_ VGND VGND VPWR VPWR _05974_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_125_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10655_ _02895_ _02925_ VGND VGND VPWR VPWR _02926_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13374_ _05366_ _05375_ VGND VGND VPWR VPWR _05899_ sky130_fd_sc_hd__nand2_1
XFILLER_0_140_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10586_ _04895_ _04928_ _02849_ _02304_ VGND VGND VPWR VPWR _02851_ sky130_fd_sc_hd__and4_1
XFILLER_0_24_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12325_ _01289_ _04748_ _04747_ VGND VGND VPWR VPWR _04762_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_51_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__07429__D _04059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12256_ _04678_ _04684_ _04685_ VGND VGND VPWR VPWR _04687_ sky130_fd_sc_hd__or3_1
XANTENNA__12632__B _00392_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11207_ _03514_ _03533_ VGND VGND VPWR VPWR _03534_ sky130_fd_sc_hd__and2b_1
XFILLER_0_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12187_ _03613_ _03623_ VGND VGND VPWR VPWR _04611_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13447__C _02735_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11371__A1 _03690_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11138_ _03453_ _03457_ VGND VGND VPWR VPWR _03458_ sky130_fd_sc_hd__or2_2
X_11069_ _03379_ _03380_ VGND VGND VPWR VPWR _03382_ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09867__A2 _01260_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07300_ _00770_ _00803_ VGND VGND VPWR VPWR _02653_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08280_ _00324_ _00326_ VGND VGND VPWR VPWR _00327_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_128_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07231_ _00967_ _01011_ VGND VGND VPWR VPWR _01897_ sky130_fd_sc_hd__or2_1
XANTENNA__11711__B _00916_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07162_ _01109_ _01131_ VGND VGND VPWR VPWR _01142_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_54_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07093_ _00377_ VGND VGND VPWR VPWR _00388_ sky130_fd_sc_hd__buf_4
XANTENNA__12851__A1_N _02857_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11362__A1 _02246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11362__B2 _02249_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09803_ _01991_ _01992_ VGND VGND VPWR VPWR _01993_ sky130_fd_sc_hd__nor2_1
X_07995_ _07005_ _07034_ _07033_ VGND VGND VPWR VPWR _00039_ sky130_fd_sc_hd__a21o_1
X_09734_ _02467_ _01060_ VGND VGND VPWR VPWR _01917_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12311__B1 _01664_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07652__A _06428_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09665_ _00843_ _00670_ _00145_ _04917_ VGND VGND VPWR VPWR _01841_ sky130_fd_sc_hd__and4_1
XANTENNA__08467__B _06873_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08530__A2 _00460_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08616_ _00692_ _00693_ VGND VGND VPWR VPWR _00695_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09596_ _00475_ net10 _01615_ _01617_ VGND VGND VPWR VPWR _01767_ sky130_fd_sc_hd__a31o_1
XTAP_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08547_ _00444_ _00449_ _00618_ VGND VGND VPWR VPWR _00619_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08478_ _00543_ VGND VGND VPWR VPWR _00544_ sky130_fd_sc_hd__buf_4
XFILLER_0_64_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_555 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07429_ _00442_ _02051_ _04037_ _04059_ VGND VGND VPWR VPWR _04070_ sky130_fd_sc_hd__and4_1
XFILLER_0_64_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11621__B _01182_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10518__A _01473_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07099__A _00442_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10440_ _02439_ _02470_ VGND VGND VPWR VPWR _02691_ sky130_fd_sc_hd__and2_1
XFILLER_0_60_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09794__A1 _06417_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10371_ _02597_ _02395_ _02599_ _02614_ VGND VGND VPWR VPWR _02615_ sky130_fd_sc_hd__or4_2
XANTENNA__09794__B2 _06439_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12110_ _04429_ _04505_ _04508_ VGND VGND VPWR VPWR _04526_ sky130_fd_sc_hd__or3_1
X_13090_ _05525_ _05595_ _05603_ VGND VGND VPWR VPWR _05604_ sky130_fd_sc_hd__a21oi_1
X_12041_ _04407_ _04448_ _04406_ VGND VGND VPWR VPWR _04450_ sky130_fd_sc_hd__a21o_1
XANTENNA__11349__A _02249_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13992_ _06577_ VGND VGND VPWR VPWR _06578_ sky130_fd_sc_hd__inv_2
X_12943_ _05436_ _05439_ _05441_ VGND VGND VPWR VPWR _05442_ sky130_fd_sc_hd__and3_2
XANTENNA__08521__A2 _00389_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12874_ _05238_ _05364_ _05365_ VGND VGND VPWR VPWR _05366_ sky130_fd_sc_hd__a21o_1
XTAP_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11825_ _04193_ _04211_ VGND VGND VPWR VPWR _04212_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output102_A net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12908__A _04714_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11756_ _04135_ _02643_ _02639_ VGND VGND VPWR VPWR _04137_ sky130_fd_sc_hd__a21o_1
XFILLER_0_28_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12627__B _01060_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10707_ _02975_ _02980_ _02983_ VGND VGND VPWR VPWR _02984_ sky130_fd_sc_hd__or3_1
XFILLER_0_83_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11687_ _04054_ _04060_ VGND VGND VPWR VPWR _04061_ sky130_fd_sc_hd__xor2_1
XFILLER_0_36_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13426_ _05954_ _05955_ VGND VGND VPWR VPWR _05957_ sky130_fd_sc_hd__and2b_1
XANTENNA__09234__B1 _01369_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09001__B _01039_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10638_ _00859_ _02858_ _02907_ VGND VGND VPWR VPWR _02908_ sky130_fd_sc_hd__and3_1
XFILLER_0_125_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10919__A1 _02171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10147__B _04048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10919__B2 _02467_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13357_ _05869_ _05351_ _05878_ VGND VGND VPWR VPWR _05881_ sky130_fd_sc_hd__a21oi_1
X_10569_ _00819_ _01934_ _02831_ _02815_ VGND VGND VPWR VPWR _02832_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_11_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12308_ _04737_ _04739_ _04743_ VGND VGND VPWR VPWR _04744_ sky130_fd_sc_hd__o21a_1
XFILLER_0_11_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13288_ _05602_ _05733_ _05737_ VGND VGND VPWR VPWR _05811_ sky130_fd_sc_hd__o21a_1
XFILLER_0_20_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12239_ _04666_ _04667_ VGND VGND VPWR VPWR _04668_ sky130_fd_sc_hd__xnor2_2
XANTENNA__09952__A net52 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07780_ _05060_ _06908_ VGND VGND VPWR VPWR _06909_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput4 a[12] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_36_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09450_ _01605_ _01606_ VGND VGND VPWR VPWR _01607_ sky130_fd_sc_hd__or2_2
X_08401_ _00458_ VGND VGND VPWR VPWR _00459_ sky130_fd_sc_hd__buf_4
X_09381_ _01508_ _01399_ VGND VGND VPWR VPWR _01531_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08332_ _00383_ VGND VGND VPWR VPWR _00384_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08263_ _02040_ _00143_ _00140_ _00139_ _04917_ VGND VGND VPWR VPWR _00308_ sky130_fd_sc_hd__a32o_1
XFILLER_0_6_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07214_ _01602_ _01591_ VGND VGND VPWR VPWR _01711_ sky130_fd_sc_hd__and2b_1
X_08194_ _00234_ _00236_ _00237_ VGND VGND VPWR VPWR _00238_ sky130_fd_sc_hd__and3_1
XFILLER_0_6_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07145_ _00934_ _00945_ VGND VGND VPWR VPWR _00956_ sky130_fd_sc_hd__and2b_1
XFILLER_0_131_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09846__B _02039_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12780__B1 _02305_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__07647__A _06439_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10504__C _02720_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10801__A _06483_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07978_ _00541_ _06818_ _06821_ net30 VGND VGND VPWR VPWR _00022_ sky130_fd_sc_hd__a22o_1
XANTENNA__08478__A _00543_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07382__A _03543_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09717_ _01891_ _01898_ VGND VGND VPWR VPWR _01899_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11099__B1 _03414_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09648_ _01614_ _01621_ _01823_ VGND VGND VPWR VPWR _01824_ sky130_fd_sc_hd__a21o_2
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09579_ _01737_ _01747_ VGND VGND VPWR VPWR _01748_ sky130_fd_sc_hd__xor2_1
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11610_ _03935_ _03934_ VGND VGND VPWR VPWR _03976_ sky130_fd_sc_hd__xnor2_1
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12590_ _00915_ _00916_ _02855_ _02857_ VGND VGND VPWR VPWR _05054_ sky130_fd_sc_hd__nand4_2
XFILLER_0_92_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11541_ _06873_ _01247_ _01564_ _06874_ VGND VGND VPWR VPWR _03900_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09459__D net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11472_ _03801_ _03803_ _03807_ VGND VGND VPWR VPWR _03824_ sky130_fd_sc_hd__or3_1
XANTENNA__08941__A _00943_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13211_ _05734_ _05735_ _05736_ VGND VGND VPWR VPWR _05737_ sky130_fd_sc_hd__a21o_1
X_10423_ _00311_ net24 _02460_ _02462_ VGND VGND VPWR VPWR _02672_ sky130_fd_sc_hd__a31o_1
X_14191_ _06635_ _06697_ VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__xor2_4
XFILLER_0_33_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07557__A _05467_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13142_ _05637_ _05638_ VGND VGND VPWR VPWR _05661_ sky130_fd_sc_hd__xnor2_2
X_10354_ _02594_ _02436_ _02595_ VGND VGND VPWR VPWR _02596_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_131_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13073_ _02709_ _02710_ _05584_ VGND VGND VPWR VPWR _05585_ sky130_fd_sc_hd__and3_1
XFILLER_0_130_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10285_ _02159_ _02505_ _02506_ _02519_ VGND VGND VPWR VPWR _02520_ sky130_fd_sc_hd__and4_1
X_12024_ _04429_ _04430_ VGND VGND VPWR VPWR _04431_ sky130_fd_sc_hd__nor2_1
XANTENNA__09772__A _00344_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09491__B _04169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08388__A _00978_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07292__A net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13975_ _06553_ _06555_ VGND VGND VPWR VPWR _06559_ sky130_fd_sc_hd__nand2_1
XANTENNA__07723__C _03510_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12926_ _05421_ _05422_ VGND VGND VPWR VPWR _05424_ sky130_fd_sc_hd__nand2b_2
XTAP_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13741__B _02855_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12857_ _05341_ _05347_ VGND VGND VPWR VPWR _05348_ sky130_fd_sc_hd__xor2_1
XTAP_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_831 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11808_ _04151_ _04156_ _04163_ VGND VGND VPWR VPWR _04194_ sky130_fd_sc_hd__and3_1
XFILLER_0_28_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12788_ _05266_ _05271_ VGND VGND VPWR VPWR _05272_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_145_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11899__D _03682_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11739_ _00654_ _01188_ _01289_ _00543_ VGND VGND VPWR VPWR _04118_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_28_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08851__A _03268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13409_ _05248_ _05400_ _05399_ VGND VGND VPWR VPWR _05938_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10605__B _01412_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08950_ _01058_ VGND VGND VPWR VPWR _01059_ sky130_fd_sc_hd__clkbuf_4
X_07901_ _07018_ _07029_ VGND VGND VPWR VPWR _07030_ sky130_fd_sc_hd__nor2_1
X_08881_ _00981_ _00983_ VGND VGND VPWR VPWR _00984_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_138_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07832_ _06870_ _06960_ VGND VGND VPWR VPWR _06961_ sky130_fd_sc_hd__nor2_1
X_07763_ _06854_ _06891_ VGND VGND VPWR VPWR _06892_ sky130_fd_sc_hd__xnor2_1
X_09502_ _01661_ _01662_ VGND VGND VPWR VPWR _01663_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13490__A1 _01062_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07694_ _01076_ _06818_ _06820_ _01120_ VGND VGND VPWR VPWR _06823_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09433_ _00157_ _01585_ _01587_ _01276_ VGND VGND VPWR VPWR _01588_ sky130_fd_sc_hd__nand4_1
XFILLER_0_94_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09364_ _01375_ _01378_ _01511_ VGND VGND VPWR VPWR _01512_ sky130_fd_sc_hd__o21a_1
XFILLER_0_59_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08315_ _00089_ _00184_ _00090_ VGND VGND VPWR VPWR _00365_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_129_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09295_ _00898_ _01434_ _01436_ VGND VGND VPWR VPWR _01437_ sky130_fd_sc_hd__o21bai_4
XFILLER_0_7_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10068__A _02246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08246_ _00287_ _00289_ VGND VGND VPWR VPWR _00290_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_145_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08177_ _04774_ _00220_ VGND VGND VPWR VPWR _00221_ sky130_fd_sc_hd__nor2_1
XFILLER_0_70_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07128_ _00748_ _00759_ VGND VGND VPWR VPWR _00770_ sky130_fd_sc_hd__xnor2_2
XANTENNA__07377__A net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10764__C1 _02766_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10070_ _02253_ _02283_ VGND VGND VPWR VPWR _02285_ sky130_fd_sc_hd__nor2_1
X_13760_ _06320_ _06322_ VGND VGND VPWR VPWR _06323_ sky130_fd_sc_hd__nand2_1
X_10972_ _00145_ _00460_ _03272_ _03273_ VGND VGND VPWR VPWR _03275_ sky130_fd_sc_hd__a22oi_1
XANTENNA__12284__A2 _01182_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12711_ _00393_ _01062_ _01415_ _00391_ VGND VGND VPWR VPWR _05187_ sky130_fd_sc_hd__a22o_1
X_13691_ _02088_ _02720_ _06246_ VGND VGND VPWR VPWR _06247_ sky130_fd_sc_hd__and3_1
XFILLER_0_78_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12642_ _05056_ _05110_ VGND VGND VPWR VPWR _05111_ sky130_fd_sc_hd__xor2_2
XFILLER_0_38_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13233__A1 _02278_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12573_ _04898_ _04909_ _04926_ _05033_ _05034_ VGND VGND VPWR VPWR _05035_ sky130_fd_sc_hd__a221o_1
XANTENNA__09189__D _00818_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07999__B1 _04939_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11524_ _03863_ _03864_ VGND VGND VPWR VPWR _03881_ sky130_fd_sc_hd__nor2_1
XANTENNA__09767__A _01953_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13289__A _05789_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11455_ _03543_ _02673_ VGND VGND VPWR VPWR _03805_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12624__C _02849_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10406_ _02029_ _01564_ _02448_ _02450_ VGND VGND VPWR VPWR _02654_ sky130_fd_sc_hd__a31o_1
X_14174_ _06772_ _06773_ _06636_ _06752_ _06759_ VGND VGND VPWR VPWR _06774_ sky130_fd_sc_hd__a2111o_1
XANTENNA__08412__A1 _02149_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11386_ _03724_ _03727_ VGND VGND VPWR VPWR _03730_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08412__B2 _05588_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10425__B _02673_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13439__D _02726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13125_ _05637_ _05638_ VGND VGND VPWR VPWR _05642_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10337_ _02563_ _02577_ VGND VGND VPWR VPWR _02578_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_103_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10144__C _04015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13056_ _02592_ _02703_ _02593_ VGND VGND VPWR VPWR _05567_ sky130_fd_sc_hd__a21boi_2
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10268_ _02500_ _02344_ _02501_ VGND VGND VPWR VPWR _02502_ sky130_fd_sc_hd__o21ai_4
XANTENNA__12640__B _02855_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12007_ _04329_ _04333_ _04412_ VGND VGND VPWR VPWR _04413_ sky130_fd_sc_hd__o21a_1
XANTENNA__09912__A1 _03070_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09912__B2 _02335_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10199_ _02090_ VGND VGND VPWR VPWR _02427_ sky130_fd_sc_hd__clkbuf_4
X_13958_ _06537_ _06540_ VGND VGND VPWR VPWR _06541_ sky130_fd_sc_hd__or2_1
XANTENNA__07172__D _00573_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12909_ _05403_ _05404_ VGND VGND VPWR VPWR _05405_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13889_ _06457_ _06460_ _06463_ _06464_ VGND VGND VPWR VPWR _06465_ sky130_fd_sc_hd__a211o_1
XANTENNA__08565__B _00508_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_706 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09979__A1 _06637_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11235__B1 _01415_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_683 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08100_ _00143_ VGND VGND VPWR VPWR _00144_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__10589__A2 _01413_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09080_ _00929_ _01201_ VGND VGND VPWR VPWR _01202_ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08581__A _00388_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08651__B2 _01470_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08031_ _00046_ _00074_ VGND VGND VPWR VPWR _00075_ sky130_fd_sc_hd__xor2_2
Xinput40 b[16] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__buf_4
XANTENNA__10038__D _02247_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_142_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput51 b[26] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__clkbuf_2
Xinput62 b[7] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_12_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13349__D _02857_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09982_ _01505_ VGND VGND VPWR VPWR _02189_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_110_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07347__D net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08933_ _01034_ _01040_ VGND VGND VPWR VPWR _01041_ sky130_fd_sc_hd__xor2_2
XFILLER_0_42_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08706__A2 net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08864_ _01230_ net45 VGND VGND VPWR VPWR _00965_ sky130_fd_sc_hd__and2_1
XANTENNA__10351__A _02496_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07815_ _06942_ _06943_ VGND VGND VPWR VPWR _06944_ sky130_fd_sc_hd__xnor2_1
X_08795_ _00631_ _00715_ _00598_ VGND VGND VPWR VPWR _00890_ sky130_fd_sc_hd__o21bai_1
X_07746_ _06874_ VGND VGND VPWR VPWR _06875_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__13463__A1 _01252_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07677_ _06744_ VGND VGND VPWR VPWR _06775_ sky130_fd_sc_hd__buf_4
XFILLER_0_67_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09416_ _01567_ _01564_ _00311_ _01565_ VGND VGND VPWR VPWR _01570_ sky130_fd_sc_hd__and4b_1
XANTENNA__08890__A1 _06966_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08890__B2 _06965_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09347_ _02960_ _04015_ _04180_ _00355_ VGND VGND VPWR VPWR _01494_ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11777__A1 _05456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11777__B2 _05478_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09278_ _01058_ _01418_ VGND VGND VPWR VPWR _01419_ sky130_fd_sc_hd__and2_1
XFILLER_0_133_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08229_ _00271_ _00272_ VGND VGND VPWR VPWR _00273_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_90_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11240_ _03221_ _03239_ VGND VGND VPWR VPWR _03570_ sky130_fd_sc_hd__xor2_2
XFILLER_0_105_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11171_ _03053_ _03493_ VGND VGND VPWR VPWR _03494_ sky130_fd_sc_hd__or2_1
XFILLER_0_101_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12741__A _00783_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10122_ _02340_ _02341_ VGND VGND VPWR VPWR _02342_ sky130_fd_sc_hd__nor2_2
XANTENNA__07835__A _06873_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10053_ _01859_ _01865_ _02265_ VGND VGND VPWR VPWR _02267_ sky130_fd_sc_hd__or3b_1
XFILLER_0_100_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13812_ _06377_ _06379_ VGND VGND VPWR VPWR _06380_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10955_ _04895_ _01507_ _01504_ _04928_ VGND VGND VPWR VPWR _03256_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13743_ _06301_ _06303_ VGND VGND VPWR VPWR _06304_ sky130_fd_sc_hd__xor2_1
XANTENNA__08330__B1 _00381_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12619__C _01060_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13674_ _06214_ _06227_ VGND VGND VPWR VPWR _06228_ sky130_fd_sc_hd__xor2_2
XFILLER_0_39_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07684__A2 net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10886_ _03166_ _03179_ VGND VGND VPWR VPWR _03181_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12625_ _00572_ _01411_ _02306_ _00414_ VGND VGND VPWR VPWR _05092_ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09497__A _04268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12556_ _05000_ _05015_ VGND VGND VPWR VPWR _05017_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_136_571 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12635__B _01933_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11507_ _03781_ _03780_ VGND VGND VPWR VPWR _03863_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12487_ _04937_ _04938_ _04940_ VGND VGND VPWR VPWR _04941_ sky130_fd_sc_hd__and3_1
XFILLER_0_110_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11438_ _00843_ _03783_ _03786_ VGND VGND VPWR VPWR _03787_ sky130_fd_sc_hd__and3_1
X_14226_ _00224_ _00231_ VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__xor2_2
XANTENNA_output94_A net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10155__B _02377_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_427 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13390__B1 _02673_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14157_ _05959_ _06753_ VGND VGND VPWR VPWR _06757_ sky130_fd_sc_hd__or2_1
X_11369_ _03692_ net142 _03710_ VGND VGND VPWR VPWR _03711_ sky130_fd_sc_hd__o21a_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07745__A _06821_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13108_ _05605_ _05623_ VGND VGND VPWR VPWR _05624_ sky130_fd_sc_hd__nor2_1
X_14088_ _06681_ _06682_ VGND VGND VPWR VPWR _06683_ sky130_fd_sc_hd__xnor2_4
XANTENNA__13466__B _02722_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13039_ _05541_ _05547_ VGND VGND VPWR VPWR _05548_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_119_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10602__C _00142_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07372__A1 _02456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07600_ _05808_ _05923_ VGND VGND VPWR VPWR _05934_ sky130_fd_sc_hd__nor2_1
X_08580_ _00399_ _00654_ _00543_ _03015_ VGND VGND VPWR VPWR _00655_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07531_ _04378_ VGND VGND VPWR VPWR _05192_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_49_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08295__B _00342_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07462_ net58 net32 net2 net163 VGND VGND VPWR VPWR _04433_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_847 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09201_ _06965_ _06966_ _00143_ _00158_ VGND VGND VPWR VPWR _01334_ sky130_fd_sc_hd__and4_1
XFILLER_0_119_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07393_ _03664_ VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_146_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09132_ _01193_ _01199_ VGND VGND VPWR VPWR _01258_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_856 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09063_ _01182_ VGND VGND VPWR VPWR _01183_ sky130_fd_sc_hd__buf_4
XFILLER_0_72_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09557__D _07040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08014_ _07058_ _07063_ VGND VGND VPWR VPWR _00058_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12561__A _00390_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09965_ _02051_ _01934_ _02169_ _00453_ VGND VGND VPWR VPWR _02170_ sky130_fd_sc_hd__a22o_1
XANTENNA__10081__A _02293_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08916_ _00817_ _00821_ _01021_ _00645_ VGND VGND VPWR VPWR _01023_ sky130_fd_sc_hd__a211oi_2
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09896_ _02089_ _02093_ VGND VGND VPWR VPWR _02095_ sky130_fd_sc_hd__and2_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10512__C _02765_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08847_ _00944_ _00946_ VGND VGND VPWR VPWR _00947_ sky130_fd_sc_hd__or2b_1
XANTENNA__10231__D net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08778_ _00857_ _00871_ VGND VGND VPWR VPWR _00872_ sky130_fd_sc_hd__xnor2_2
XANTENNA__13436__A1 _05833_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07729_ net28 net64 _06820_ _00563_ VGND VGND VPWR VPWR _06858_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10740_ _02987_ _03019_ VGND VGND VPWR VPWR _03020_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__08863__A1 _01284_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10671_ _05181_ _02849_ _02304_ _00094_ VGND VGND VPWR VPWR _02944_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12410_ _04854_ _04855_ VGND VGND VPWR VPWR _04856_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_63_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13390_ _00779_ _03681_ _02673_ _01518_ VGND VGND VPWR VPWR _05917_ sky130_fd_sc_hd__a22o_1
X_12341_ _03729_ _03762_ _01368_ _00959_ VGND VGND VPWR VPWR _04780_ sky130_fd_sc_hd__and4_1
XFILLER_0_106_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12272_ _04673_ _04703_ VGND VGND VPWR VPWR _04704_ sky130_fd_sc_hd__xnor2_1
X_14011_ _06509_ _06519_ _06518_ VGND VGND VPWR VPWR _06599_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_105_298 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11223_ _03548_ _03549_ _03550_ VGND VGND VPWR VPWR _03551_ sky130_fd_sc_hd__a21o_1
XFILLER_0_31_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09040__A1 _01155_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07565__A _03268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13286__B _05807_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11154_ _03473_ _03474_ VGND VGND VPWR VPWR _03475_ sky130_fd_sc_hd__xnor2_2
XANTENNA__10703__B _03004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10105_ _00628_ _05742_ net50 _01545_ VGND VGND VPWR VPWR _02323_ sky130_fd_sc_hd__and4_1
XANTENNA__07284__B _02467_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11085_ _03394_ _03395_ VGND VGND VPWR VPWR _03399_ sky130_fd_sc_hd__and2_1
X_10036_ _00844_ VGND VGND VPWR VPWR _02249_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_86_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11987_ _04287_ _04321_ VGND VGND VPWR VPWR _04391_ sky130_fd_sc_hd__and2b_1
XFILLER_0_105_24 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13726_ _06259_ _06261_ VGND VGND VPWR VPWR _06286_ sky130_fd_sc_hd__xnor2_1
X_10938_ _03231_ _03223_ VGND VGND VPWR VPWR _03238_ sky130_fd_sc_hd__and2b_1
XFILLER_0_105_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13657_ _06165_ _06163_ VGND VGND VPWR VPWR _06210_ sky130_fd_sc_hd__and2b_1
X_10869_ _03149_ _03152_ _03153_ VGND VGND VPWR VPWR _03162_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_38_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12608_ _05063_ _05062_ VGND VGND VPWR VPWR _05074_ sky130_fd_sc_hd__and2b_1
XPHY_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13588_ _01414_ _03783_ _06124_ VGND VGND VPWR VPWR _06134_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_143_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09020__A _06966_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12539_ _04817_ _04997_ VGND VGND VPWR VPWR _04998_ sky130_fd_sc_hd__nand2_2
XFILLER_0_30_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09955__A _04081_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07290__B1 net61 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14209_ _01733_ _01755_ VGND VGND VPWR VPWR _06799_ sky130_fd_sc_hd__or2_1
XFILLER_0_112_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09750_ _00453_ _01934_ VGND VGND VPWR VPWR _01935_ sky130_fd_sc_hd__and2_1
X_08701_ _00776_ _00786_ VGND VGND VPWR VPWR _00787_ sky130_fd_sc_hd__xor2_2
XANTENNA__09690__A _04939_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09681_ _01857_ _01858_ VGND VGND VPWR VPWR _01859_ sky130_fd_sc_hd__and2_1
XANTENNA__11677__B1 _01260_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08632_ _00551_ _00347_ _00711_ VGND VGND VPWR VPWR _00712_ sky130_fd_sc_hd__and3b_1
XFILLER_0_146_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08563_ _00635_ VGND VGND VPWR VPWR _00636_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_89_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07514_ net44 _04851_ net4 _00573_ VGND VGND VPWR VPWR _05005_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_222 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08494_ _00559_ _00560_ VGND VGND VPWR VPWR _00561_ sky130_fd_sc_hd__and2b_1
XFILLER_0_77_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07445_ _04224_ _04235_ VGND VGND VPWR VPWR _04246_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_64_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07376_ _02894_ _03477_ VGND VGND VPWR VPWR _03488_ sky130_fd_sc_hd__xor2_4
XFILLER_0_18_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09115_ _00727_ _00893_ _00899_ VGND VGND VPWR VPWR _01240_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_72_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10955__A2 _01507_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09046_ _01163_ VGND VGND VPWR VPWR _01165_ sky130_fd_sc_hd__inv_2
XANTENNA__09865__A _06765_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13818__C _03686_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07385__A _00978_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09948_ _01942_ _01944_ VGND VGND VPWR VPWR _02152_ sky130_fd_sc_hd__nor2_1
X_09879_ _02074_ _02075_ VGND VGND VPWR VPWR _02076_ sky130_fd_sc_hd__nand2_1
X_11910_ _04201_ _04210_ VGND VGND VPWR VPWR _04306_ sky130_fd_sc_hd__nand2_1
XTAP_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12890_ _01954_ _05220_ _05222_ _05223_ VGND VGND VPWR VPWR _05384_ sky130_fd_sc_hd__o2bb2ai_1
XTAP_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09105__A _00530_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11841_ _04223_ _04226_ VGND VGND VPWR VPWR _04230_ sky130_fd_sc_hd__nand2_1
XTAP_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_542 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11772_ _04152_ _04153_ _01996_ net20 VGND VGND VPWR VPWR _04154_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_68_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13511_ _05985_ _02722_ _05998_ _05997_ VGND VGND VPWR VPWR _06049_ sky130_fd_sc_hd__a31o_1
X_10723_ _02998_ _03000_ VGND VGND VPWR VPWR _03001_ sky130_fd_sc_hd__or2_2
XTAP_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10654_ _02842_ _02893_ VGND VGND VPWR VPWR _02925_ sky130_fd_sc_hd__or2_1
X_13442_ _05969_ _02765_ _05971_ _05972_ VGND VGND VPWR VPWR _05973_ sky130_fd_sc_hd__and4_1
XFILLER_0_137_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12396__A1 _00374_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13373_ _05896_ _05897_ VGND VGND VPWR VPWR _05898_ sky130_fd_sc_hd__and2_1
X_10585_ _02158_ VGND VGND VPWR VPWR _02849_ sky130_fd_sc_hd__buf_2
XFILLER_0_134_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12324_ _04759_ _04760_ VGND VGND VPWR VPWR _04761_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12255_ _04665_ _04668_ VGND VGND VPWR VPWR _04685_ sky130_fd_sc_hd__xor2_1
XFILLER_0_121_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11206_ _03518_ _03530_ _03531_ VGND VGND VPWR VPWR _03533_ sky130_fd_sc_hd__o21ba_1
XANTENNA__12632__C _02723_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12186_ _04602_ _04606_ _04607_ _04608_ VGND VGND VPWR VPWR _04610_ sky130_fd_sc_hd__a211o_1
XANTENNA__13447__D _02731_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11137_ _03450_ _03452_ VGND VGND VPWR VPWR _03457_ sky130_fd_sc_hd__nor2_1
X_11068_ _03379_ _03380_ VGND VGND VPWR VPWR _03381_ sky130_fd_sc_hd__nand2_1
XANTENNA__07327__A1 _00344_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10019_ _04862_ _04873_ _04037_ _04059_ VGND VGND VPWR VPWR _02230_ sky130_fd_sc_hd__and4_1
XFILLER_0_58_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08827__A1 _00901_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13820__A1 _01955_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_575 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13709_ _06265_ _06266_ VGND VGND VPWR VPWR _06267_ sky130_fd_sc_hd__xor2_1
XFILLER_0_86_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07230_ _00858_ _01875_ VGND VGND VPWR VPWR _01886_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_144_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12387__A1 _00374_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07161_ _01120_ net59 VGND VGND VPWR VPWR _01131_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07092_ _00366_ VGND VGND VPWR VPWR _00377_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_112_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11898__B1 _02135_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11362__A2 _03687_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09802_ _01782_ _01784_ _01990_ VGND VGND VPWR VPWR _01992_ sky130_fd_sc_hd__nor3_1
X_07994_ _00007_ _00037_ VGND VGND VPWR VPWR _00038_ sky130_fd_sc_hd__xor2_1
X_09733_ _01912_ _01915_ VGND VGND VPWR VPWR _01916_ sky130_fd_sc_hd__xor2_2
XANTENNA__12311__A1 _00607_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12311__B2 _00415_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11455__A _03543_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07652__B _06450_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09664_ _00843_ _00635_ _01839_ VGND VGND VPWR VPWR _01840_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_69_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08467__C _06875_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08615_ _00500_ _00502_ _00691_ VGND VGND VPWR VPWR _00693_ sky130_fd_sc_hd__nor3_1
X_09595_ _01763_ _01764_ VGND VGND VPWR VPWR _01765_ sky130_fd_sc_hd__xor2_1
XTAP_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13670__A _01183_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08546_ _00611_ _00616_ VGND VGND VPWR VPWR _00618_ sky130_fd_sc_hd__xor2_1
X_08477_ _07004_ VGND VGND VPWR VPWR _00543_ sky130_fd_sc_hd__buf_4
XFILLER_0_65_748 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07428_ _04048_ VGND VGND VPWR VPWR _04059_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_92_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_636 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10518__B _02722_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07359_ _01295_ _01405_ _02664_ _02719_ VGND VGND VPWR VPWR _03301_ sky130_fd_sc_hd__nand4_2
XFILLER_0_45_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10370_ _02612_ _02613_ VGND VGND VPWR VPWR _02614_ sky130_fd_sc_hd__nor2_1
XANTENNA__09794__A2 _00574_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09029_ _01144_ _01145_ VGND VGND VPWR VPWR _01146_ sky130_fd_sc_hd__and2_1
XFILLER_0_103_544 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12040_ _04407_ _04448_ VGND VGND VPWR VPWR _04449_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11349__B _01312_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_split3_A _00869_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08939__A _00991_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13991_ _06568_ _06574_ _06576_ VGND VGND VPWR VPWR _06577_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_99_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12942_ _02391_ _02150_ _02479_ _05440_ _05438_ VGND VGND VPWR VPWR _05441_ sky130_fd_sc_hd__a2111o_2
XTAP_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12873_ _00458_ _03748_ _05239_ VGND VGND VPWR VPWR _05365_ sky130_fd_sc_hd__and3_1
XTAP_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13580__A _01414_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11824_ _04201_ _04210_ VGND VGND VPWR VPWR _04211_ sky130_fd_sc_hd__xnor2_1
XTAP_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12908__B _01957_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10616__A1 _01472_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11755_ _02634_ _02637_ VGND VGND VPWR VPWR _04135_ sky130_fd_sc_hd__or2b_1
XFILLER_0_55_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10706_ _02970_ _02981_ VGND VGND VPWR VPWR _02983_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11686_ _02407_ _02611_ _04057_ _04058_ VGND VGND VPWR VPWR _04060_ sky130_fd_sc_hd__o31a_1
X_13425_ _05413_ _05852_ _05953_ VGND VGND VPWR VPWR _05955_ sky130_fd_sc_hd__a21o_1
XANTENNA__09234__A1 _04268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10637_ _01472_ _02856_ VGND VGND VPWR VPWR _02907_ sky130_fd_sc_hd__nand2_1
XFILLER_0_141_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09234__B2 _01372_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10919__A2 _02758_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10147__C _05027_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10568_ _02814_ VGND VGND VPWR VPWR _02831_ sky130_fd_sc_hd__inv_2
X_13356_ _05869_ _05351_ _05878_ VGND VGND VPWR VPWR _05880_ sky130_fd_sc_hd__and3_1
XFILLER_0_106_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12307_ _04740_ _04742_ VGND VGND VPWR VPWR _04743_ sky130_fd_sc_hd__xnor2_1
X_13287_ _05762_ _05764_ _05765_ _05809_ VGND VGND VPWR VPWR _05810_ sky130_fd_sc_hd__a31o_2
X_10499_ _02738_ _02739_ _02734_ VGND VGND VPWR VPWR _02755_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_121_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12362__C net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11259__B _03571_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12238_ _00375_ _02120_ VGND VGND VPWR VPWR _04667_ sky130_fd_sc_hd__nand2_1
X_12169_ _04588_ _04589_ _04590_ VGND VGND VPWR VPWR _04591_ sky130_fd_sc_hd__o21bai_1
Xinput5 a[13] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_127_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08400_ _00457_ VGND VGND VPWR VPWR _00458_ sky130_fd_sc_hd__clkbuf_4
X_09380_ _02160_ _00605_ _01508_ _02116_ VGND VGND VPWR VPWR _01530_ sky130_fd_sc_hd__a22o_1
XANTENNA__13501__A2_N _03680_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08331_ _04070_ _00382_ VGND VGND VPWR VPWR _00383_ sky130_fd_sc_hd__or2_1
XFILLER_0_52_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08262_ _03059_ _00144_ _00304_ _00305_ VGND VGND VPWR VPWR _00307_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_144_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07213_ _01624_ _01678_ _01689_ VGND VGND VPWR VPWR _01700_ sky130_fd_sc_hd__nand3_2
XFILLER_0_27_472 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08193_ _00210_ _00214_ _00208_ VGND VGND VPWR VPWR _00237_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_144_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07144_ _00420_ net61 net60 net176 VGND VGND VPWR VPWR _00945_ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_691 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_604 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12780__A1 _00572_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12780__B2 _00414_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08736__B1 _06765_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10504__D _02726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07663__A _06428_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07977_ _02719_ _03499_ _07024_ _07023_ VGND VGND VPWR VPWR _00021_ sky130_fd_sc_hd__a31o_1
XANTENNA__10801__B _01933_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09716_ _01895_ _01896_ VGND VGND VPWR VPWR _01898_ sky130_fd_sc_hd__nor2_1
XANTENNA__11099__B2 _07040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12296__B1 _02088_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09161__B1 _01289_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09647_ _01614_ _01621_ _01572_ VGND VGND VPWR VPWR _01823_ sky130_fd_sc_hd__o21a_1
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11913__A _00157_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_704 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09578_ _01745_ _01746_ VGND VGND VPWR VPWR _01747_ sky130_fd_sc_hd__nor2_1
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12599__A1 _00914_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08529_ _00454_ _00455_ _00461_ VGND VGND VPWR VPWR _00599_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_65_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13260__A2 _05779_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11540_ _06819_ _06874_ _01247_ net19 VGND VGND VPWR VPWR _03899_ sky130_fd_sc_hd__and4_1
XFILLER_0_53_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10248__B _02150_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11471_ _00519_ _03679_ _03816_ _03822_ VGND VGND VPWR VPWR _03823_ sky130_fd_sc_hd__a31o_1
XFILLER_0_123_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13210_ _05715_ _05724_ VGND VGND VPWR VPWR _05736_ sky130_fd_sc_hd__nor2_1
X_10422_ _02669_ _02670_ VGND VGND VPWR VPWR _02671_ sky130_fd_sc_hd__xor2_1
XANTENNA__07838__A _01383_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14190_ _06632_ _06689_ VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__xor2_4
XFILLER_0_116_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_637 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13141_ _05655_ _05659_ VGND VGND VPWR VPWR _05660_ sky130_fd_sc_hd__nor2_2
X_10353_ _02095_ _02429_ _02432_ _02092_ VGND VGND VPWR VPWR _02595_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_131_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10782__B1 _02730_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13072_ _02055_ _02272_ _02488_ _05583_ VGND VGND VPWR VPWR _05584_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_130_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10284_ _02517_ _02518_ VGND VGND VPWR VPWR _02519_ sky130_fd_sc_hd__nand2_1
X_12023_ _06626_ _03683_ _03679_ _06450_ VGND VGND VPWR VPWR _04430_ sky130_fd_sc_hd__a22oi_1
XANTENNA__09772__B _01958_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08669__A _05731_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09491__C net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08388__B _00880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07292__B net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13974_ _06160_ _06557_ VGND VGND VPWR VPWR _06558_ sky130_fd_sc_hd__nand2_1
XANTENNA__07723__D _00475_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12925_ _05420_ _04629_ _05316_ VGND VGND VPWR VPWR _05422_ sky130_fd_sc_hd__or3_1
XFILLER_0_88_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12856_ _05344_ _05345_ VGND VGND VPWR VPWR _05347_ sky130_fd_sc_hd__xnor2_1
XTAP_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11807_ _04171_ _04192_ VGND VGND VPWR VPWR _04193_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_843 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12787_ _05268_ _05270_ VGND VGND VPWR VPWR _05271_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_29_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11738_ _04113_ _04116_ VGND VGND VPWR VPWR _04117_ sky130_fd_sc_hd__or2_1
XFILLER_0_113_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_455 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_88 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11669_ _06733_ _03773_ _02601_ _02600_ _03696_ VGND VGND VPWR VPWR _04041_ sky130_fd_sc_hd__a32o_1
XFILLER_0_98_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08851__B net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13408_ _05931_ _05936_ VGND VGND VPWR VPWR _05937_ sky130_fd_sc_hd__xor2_2
XFILLER_0_126_499 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07748__A _01350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13339_ _05326_ _05331_ _05860_ VGND VGND VPWR VPWR _05861_ sky130_fd_sc_hd__and3_1
XFILLER_0_11_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09963__A net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07900_ _06949_ _07028_ VGND VGND VPWR VPWR _07029_ sky130_fd_sc_hd__xnor2_1
X_08880_ _00629_ _00802_ _00982_ VGND VGND VPWR VPWR _00983_ sky130_fd_sc_hd__a21o_1
XANTENNA__08579__A _00004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07483__A _00661_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07831_ _06956_ _06959_ VGND VGND VPWR VPWR _06960_ sky130_fd_sc_hd__xnor2_1
X_07762_ _06790_ _06850_ VGND VGND VPWR VPWR _06891_ sky130_fd_sc_hd__xnor2_1
X_09501_ _01552_ _01660_ VGND VGND VPWR VPWR _01662_ sky130_fd_sc_hd__nor2_1
X_07693_ _00891_ _01120_ _06819_ _06821_ VGND VGND VPWR VPWR _06822_ sky130_fd_sc_hd__nand4_1
XFILLER_0_2_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09694__A1 _04378_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09694__B2 _02971_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09432_ _00159_ _01586_ VGND VGND VPWR VPWR _01587_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09363_ _01502_ _01510_ VGND VGND VPWR VPWR _01511_ sky130_fd_sc_hd__xor2_1
XFILLER_0_19_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08314_ _00356_ _06999_ _00357_ _00363_ VGND VGND VPWR VPWR _00364_ sky130_fd_sc_hd__or4_4
XFILLER_0_47_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09294_ _01056_ _01435_ _01238_ VGND VGND VPWR VPWR _01436_ sky130_fd_sc_hd__o21a_1
XFILLER_0_90_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10068__B _02247_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08245_ _00134_ _00136_ _00288_ VGND VGND VPWR VPWR _00289_ sky130_fd_sc_hd__a21o_1
XFILLER_0_7_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08176_ _03037_ _04763_ VGND VGND VPWR VPWR _00220_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07127_ _00541_ _00661_ VGND VGND VPWR VPWR _00759_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10764__B1 _01156_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10971_ _00142_ _00457_ _03272_ _03273_ VGND VGND VPWR VPWR _03274_ sky130_fd_sc_hd__and4_1
XFILLER_0_69_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12710_ _05184_ _05185_ VGND VGND VPWR VPWR _05186_ sky130_fd_sc_hd__nor2_1
XFILLER_0_69_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13690_ _06243_ _06245_ VGND VGND VPWR VPWR _06246_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12641_ _00916_ _02857_ _05109_ VGND VGND VPWR VPWR _05110_ sky130_fd_sc_hd__and3_1
XFILLER_0_66_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12572_ _04913_ _04925_ VGND VGND VPWR VPWR _05034_ sky130_fd_sc_hd__nor2_1
XANTENNA__08952__A _01060_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07999__A1 _02335_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07999__B2 _03070_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11523_ _03878_ _03879_ VGND VGND VPWR VPWR _03880_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07568__A _01405_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13289__B _05807_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11454_ _03792_ _03791_ VGND VGND VPWR VPWR _03804_ sky130_fd_sc_hd__and2b_1
XFILLER_0_21_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10405_ _02650_ _02651_ VGND VGND VPWR VPWR _02652_ sky130_fd_sc_hd__xor2_1
X_11385_ _03724_ _03727_ VGND VGND VPWR VPWR _03728_ sky130_fd_sc_hd__and2_1
X_14173_ _06642_ _06753_ _06613_ VGND VGND VPWR VPWR _06773_ sky130_fd_sc_hd__or3b_1
XFILLER_0_33_294 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_434 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08412__A2 _00112_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13124_ _05216_ _05640_ VGND VGND VPWR VPWR _05641_ sky130_fd_sc_hd__nand2_2
XFILLER_0_131_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10336_ _02574_ _02575_ VGND VGND VPWR VPWR _02577_ sky130_fd_sc_hd__nand2_2
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11818__A _00159_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13055_ _05556_ _05564_ VGND VGND VPWR VPWR _05565_ sky130_fd_sc_hd__nor2_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10267_ _02195_ _02338_ _02341_ _02192_ VGND VGND VPWR VPWR _02501_ sky130_fd_sc_hd__a211oi_2
XANTENNA__08399__A net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12006_ _04409_ _04410_ VGND VGND VPWR VPWR _04412_ sky130_fd_sc_hd__nor2_1
XANTENNA__09912__A2 _01180_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10198_ _02088_ VGND VGND VPWR VPWR _02426_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13957_ _06476_ _06539_ VGND VGND VPWR VPWR _06540_ sky130_fd_sc_hd__xnor2_2
XANTENNA__12649__A _02008_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12908_ _04714_ _01957_ VGND VGND VPWR VPWR _05404_ sky130_fd_sc_hd__nand2_1
X_13888_ _06462_ _06449_ VGND VGND VPWR VPWR _06464_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08565__C _04917_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12839_ _00392_ _00742_ _02723_ _02727_ VGND VGND VPWR VPWR _05328_ sky130_fd_sc_hd__and4_1
XTAP_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10169__A _06965_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_567 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11235__A1 _03015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09979__A2 _01400_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11235__B2 _00410_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08651__A2 net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08581__B _02993_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08030_ _00072_ _00073_ VGND VGND VPWR VPWR _00074_ sky130_fd_sc_hd__nand2_1
XFILLER_0_114_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput30 a[7] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__buf_2
XFILLER_0_140_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput41 b[17] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__buf_1
XFILLER_0_4_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput52 b[27] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__buf_4
XFILLER_0_12_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput63 b[8] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_24_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09981_ _02187_ VGND VGND VPWR VPWR _02188_ sky130_fd_sc_hd__clkbuf_4
X_08932_ _01036_ _01039_ VGND VGND VPWR VPWR _01040_ sky130_fd_sc_hd__xor2_2
X_08863_ _01284_ net45 _00793_ _00791_ VGND VGND VPWR VPWR _00964_ sky130_fd_sc_hd__a31o_1
XANTENNA__10351__B _02498_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08102__A _02280_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07814_ _00541_ _03499_ VGND VGND VPWR VPWR _06943_ sky130_fd_sc_hd__nand2_1
X_08794_ _00765_ _00888_ VGND VGND VPWR VPWR _00889_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_79_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07745_ _06821_ VGND VGND VPWR VPWR _06874_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__13463__A2 _02737_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07678__B1 _06775_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07676_ _06733_ VGND VGND VPWR VPWR _06765_ sky130_fd_sc_hd__buf_4
X_09415_ _00322_ _01564_ _01566_ _01567_ VGND VGND VPWR VPWR _01568_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_137_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08890__A2 _04906_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09346_ _01409_ _01420_ _01491_ VGND VGND VPWR VPWR _01493_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_63_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11777__A2 _02117_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09277_ _00431_ _04169_ net50 VGND VGND VPWR VPWR _01418_ sky130_fd_sc_hd__and3_1
XFILLER_0_7_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08228_ _06461_ _00003_ VGND VGND VPWR VPWR _00272_ sky130_fd_sc_hd__nand2_1
XFILLER_0_117_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08159_ _06986_ _06987_ _06997_ VGND VGND VPWR VPWR _00203_ sky130_fd_sc_hd__nand3_1
XFILLER_0_120_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11170_ _03453_ _03492_ _03454_ VGND VGND VPWR VPWR _03493_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_30_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12741__B _00779_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10121_ _02336_ _02201_ _02339_ VGND VGND VPWR VPWR _02341_ sky130_fd_sc_hd__o21a_1
XFILLER_0_30_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10052_ _01859_ _01865_ _02265_ VGND VGND VPWR VPWR _02266_ sky130_fd_sc_hd__o21bai_2
XANTENNA__13853__A _01517_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13811_ _06377_ _06378_ _01400_ _03683_ VGND VGND VPWR VPWR _06379_ sky130_fd_sc_hd__and4bb_1
X_13742_ _02088_ _02858_ _06302_ VGND VGND VPWR VPWR _06303_ sky130_fd_sc_hd__and3_1
X_10954_ _03253_ _03254_ VGND VGND VPWR VPWR _03255_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_57_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08330__A1 _00464_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08330__B2 _02051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13673_ _06215_ _06212_ VGND VGND VPWR VPWR _06227_ sky130_fd_sc_hd__nand2_1
XANTENNA__12619__D _01413_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10885_ _03165_ _03154_ _03164_ VGND VGND VPWR VPWR _03179_ sky130_fd_sc_hd__nor3_1
XFILLER_0_128_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_651 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12624_ _00414_ _00572_ _02849_ VGND VGND VPWR VPWR _05091_ sky130_fd_sc_hd__and3_1
XANTENNA__09778__A _01306_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09497__B net49 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12555_ _04998_ _04999_ VGND VGND VPWR VPWR _05015_ sky130_fd_sc_hd__xor2_2
XFILLER_0_136_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_274 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11506_ _03859_ _03860_ VGND VGND VPWR VPWR _03862_ sky130_fd_sc_hd__or2_2
XFILLER_0_79_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12486_ _00779_ _00755_ _00741_ _00783_ VGND VGND VPWR VPWR _04940_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14225_ _06807_ _06808_ VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__nor2_2
X_11437_ _00844_ _03785_ VGND VGND VPWR VPWR _03786_ sky130_fd_sc_hd__nand2_1
XFILLER_0_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13390__A1 _00779_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14156_ _05830_ _05833_ _05962_ _06754_ VGND VGND VPWR VPWR _06756_ sky130_fd_sc_hd__o211ai_2
XANTENNA__13390__B2 _01518_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11368_ _03708_ _03709_ VGND VGND VPWR VPWR _03710_ sky130_fd_sc_hd__nor2_1
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13107_ _05622_ VGND VGND VPWR VPWR _05623_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10319_ _02361_ _02557_ VGND VGND VPWR VPWR _02558_ sky130_fd_sc_hd__nand2_1
X_14087_ _06116_ _06237_ _06115_ VGND VGND VPWR VPWR _06682_ sky130_fd_sc_hd__a21o_2
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11299_ _02770_ _02787_ VGND VGND VPWR VPWR _03635_ sky130_fd_sc_hd__nor2_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13038_ _05532_ _05539_ VGND VGND VPWR VPWR _05547_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_28_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10602__D _01059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08857__A _00431_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07372__A2 _02467_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07530_ _04598_ VGND VGND VPWR VPWR _05181_ sky130_fd_sc_hd__buf_4
XFILLER_0_88_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07461_ net58 net175 net32 net2 VGND VGND VPWR VPWR _04422_ sky130_fd_sc_hd__and4_1
XFILLER_0_76_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09200_ _00262_ _00144_ _00298_ _00263_ VGND VGND VPWR VPWR _01333_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_147_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07392_ _03642_ _03653_ VGND VGND VPWR VPWR _03664_ sky130_fd_sc_hd__and2_1
XFILLER_0_60_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09131_ _01192_ _01200_ VGND VGND VPWR VPWR _01257_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09062_ _01181_ VGND VGND VPWR VPWR _01182_ sky130_fd_sc_hd__buf_4
XFILLER_0_13_710 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08013_ _00055_ _00056_ VGND VGND VPWR VPWR _00057_ sky130_fd_sc_hd__xor2_1
XFILLER_0_115_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_592 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12561__B _01066_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09964_ _02168_ VGND VGND VPWR VPWR _02169_ sky130_fd_sc_hd__clkbuf_4
X_08915_ _00822_ _00823_ VGND VGND VPWR VPWR _01021_ sky130_fd_sc_hd__and2_1
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09895_ _02091_ _02092_ VGND VGND VPWR VPWR _02093_ sky130_fd_sc_hd__nor2_1
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10512__D _02722_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08846_ _05742_ _04103_ _04191_ _00563_ VGND VGND VPWR VPWR _00946_ sky130_fd_sc_hd__a22o_1
XANTENNA__08767__A _06626_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08777_ _00866_ _00870_ VGND VGND VPWR VPWR _00871_ sky130_fd_sc_hd__xnor2_4
X_07728_ _00563_ net28 net64 net34 VGND VGND VPWR VPWR _06857_ sky130_fd_sc_hd__and4_1
XFILLER_0_67_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_223 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07659_ _06560_ _06571_ VGND VGND VPWR VPWR _06582_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08863__A2 net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10670_ _00094_ _00151_ _02849_ _02304_ VGND VGND VPWR VPWR _02943_ sky130_fd_sc_hd__nand4_1
XFILLER_0_36_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09329_ _00544_ _01473_ VGND VGND VPWR VPWR _01474_ sky130_fd_sc_hd__nand2_1
XFILLER_0_106_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10537__A _03004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12340_ _03762_ _01368_ _00959_ _03729_ VGND VGND VPWR VPWR _04779_ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12271_ _04687_ _04694_ _04695_ VGND VGND VPWR VPWR _04703_ sky130_fd_sc_hd__a21oi_1
X_14010_ _06533_ _06596_ _06597_ VGND VGND VPWR VPWR _06598_ sky130_fd_sc_hd__a21oi_4
X_11222_ _02583_ _02586_ VGND VGND VPWR VPWR _03550_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09040__A2 _01156_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_595 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11153_ _03189_ _03205_ _03242_ _03187_ VGND VGND VPWR VPWR _03474_ sky130_fd_sc_hd__a31o_1
XANTENNA__10703__C _01059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10104_ _00650_ _01410_ _02158_ _02105_ VGND VGND VPWR VPWR _02322_ sky130_fd_sc_hd__a22oi_1
X_11084_ _03278_ _03397_ VGND VGND VPWR VPWR _03398_ sky130_fd_sc_hd__nand2_2
XFILLER_0_65_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10035_ _00859_ VGND VGND VPWR VPWR _02247_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__07581__A _00639_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output125_A net125 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11986_ _04357_ _04386_ _04387_ _04385_ VGND VGND VPWR VPWR _04390_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_36 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13725_ _06277_ _06283_ _06281_ VGND VGND VPWR VPWR _06284_ sky130_fd_sc_hd__o21a_1
X_10937_ _03225_ _03236_ VGND VGND VPWR VPWR _03237_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_85_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13656_ _01252_ _02766_ _06077_ _01183_ VGND VGND VPWR VPWR _06209_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10868_ _02534_ _03160_ VGND VGND VPWR VPWR _03161_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12607_ _05065_ _05070_ _05072_ VGND VGND VPWR VPWR _05073_ sky130_fd_sc_hd__nand3_1
XPHY_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13587_ _06130_ _06132_ VGND VGND VPWR VPWR _06133_ sky130_fd_sc_hd__and2b_1
XPHY_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10799_ _03083_ _03084_ VGND VGND VPWR VPWR _03085_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_81_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09020__B _00142_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12538_ _04815_ _04816_ VGND VGND VPWR VPWR _04997_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07459__C net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07290__A1 net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09955__B _01339_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07290__B2 _00869_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12469_ _04919_ _04920_ VGND VGND VPWR VPWR _04921_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14208_ _01788_ _06798_ VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__nor2_2
XFILLER_0_111_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07756__A _06775_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14139_ _06710_ _06700_ VGND VGND VPWR VPWR _06737_ sky130_fd_sc_hd__and2b_1
XFILLER_0_10_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09971__A _02105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08700_ _01350_ _00779_ _00785_ VGND VGND VPWR VPWR _00786_ sky130_fd_sc_hd__and3_2
XANTENNA__09690__B _00379_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11677__A1 _07010_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09680_ _01737_ _01746_ _01743_ VGND VGND VPWR VPWR _01858_ sky130_fd_sc_hd__o21a_1
XANTENNA__11677__B2 _00268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08631_ _00550_ VGND VGND VPWR VPWR _00711_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_540 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08562_ _04917_ VGND VGND VPWR VPWR _00635_ sky130_fd_sc_hd__buf_2
XFILLER_0_49_426 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07513_ _00573_ net44 _04851_ net4 VGND VGND VPWR VPWR _04994_ sky130_fd_sc_hd__and4_1
XANTENNA__10101__A1 _01934_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08493_ _00558_ _00463_ VGND VGND VPWR VPWR _00560_ sky130_fd_sc_hd__nand2_2
XFILLER_0_76_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_623 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07444_ _01372_ _04026_ VGND VGND VPWR VPWR _04235_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07375_ _03466_ _03455_ VGND VGND VPWR VPWR _03477_ sky130_fd_sc_hd__nor2_4
XANTENNA__10357__A _07010_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09114_ _01056_ _01238_ VGND VGND VPWR VPWR _01239_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_44_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09045_ _01113_ _01161_ _01114_ VGND VGND VPWR VPWR _01163_ sky130_fd_sc_hd__and3_1
XFILLER_0_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09865__B _06775_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09558__B1 _07040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09881__A _03521_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09947_ _02056_ _02037_ _02038_ _02148_ _02150_ VGND VGND VPWR VPWR _02151_ sky130_fd_sc_hd__o41a_4
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09878_ _02073_ _02059_ _02060_ VGND VGND VPWR VPWR _02075_ sky130_fd_sc_hd__nand3_1
XFILLER_0_99_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08829_ _00925_ _00926_ VGND VGND VPWR VPWR _00927_ sky130_fd_sc_hd__xor2_1
XTAP_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11840_ _04149_ _04228_ VGND VGND VPWR VPWR _04229_ sky130_fd_sc_hd__nor2_1
XANTENNA__09105__B _00391_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11771_ _05445_ _01246_ net19 _05467_ VGND VGND VPWR VPWR _04153_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_95_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12747__A _00379_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13510_ _06008_ _06047_ VGND VGND VPWR VPWR _06048_ sky130_fd_sc_hd__nor2_2
XFILLER_0_95_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10722_ _01156_ _02766_ _02999_ VGND VGND VPWR VPWR _03000_ sky130_fd_sc_hd__a21oi_1
XTAP_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09121__A net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13441_ _01250_ _02721_ _02735_ _01182_ VGND VGND VPWR VPWR _05972_ sky130_fd_sc_hd__a22o_1
X_10653_ _02921_ _02923_ VGND VGND VPWR VPWR _02924_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12396__A2 _01272_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13372_ _05320_ _05321_ _05359_ _05895_ VGND VGND VPWR VPWR _05897_ sky130_fd_sc_hd__a211o_1
XFILLER_0_118_391 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10584_ _04895_ _02306_ _02305_ _04928_ VGND VGND VPWR VPWR _02848_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07272__A1 _00453_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12323_ _04750_ _04756_ _04758_ VGND VGND VPWR VPWR _04760_ sky130_fd_sc_hd__or3_1
XFILLER_0_51_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12254_ _04681_ _04683_ VGND VGND VPWR VPWR _04684_ sky130_fd_sc_hd__and2b_1
XFILLER_0_31_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11205_ net178 _03529_ _03528_ VGND VGND VPWR VPWR _03531_ sky130_fd_sc_hd__o21a_1
XANTENNA__11098__A _01400_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12185_ _03614_ _03602_ VGND VGND VPWR VPWR _04608_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11136_ _03053_ _03454_ VGND VGND VPWR VPWR _03456_ sky130_fd_sc_hd__nor2_1
XANTENNA__10221__A2_N _01564_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11067_ _03335_ _03364_ VGND VGND VPWR VPWR _03380_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07327__A2 _00410_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10018_ _04939_ _00376_ _00379_ _04917_ VGND VGND VPWR VPWR _02229_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_59_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_746 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11969_ _04369_ _04303_ _04370_ VGND VGND VPWR VPWR _04371_ sky130_fd_sc_hd__or3_1
XANTENNA__08827__A2 _03762_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13708_ _02427_ _02759_ VGND VGND VPWR VPWR _06266_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13639_ _06169_ _06170_ VGND VGND VPWR VPWR _06190_ sky130_fd_sc_hd__nand2_1
XANTENNA__10177__A _00101_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07160_ net26 VGND VGND VPWR VPWR _01120_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__12387__A2 _01584_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09966__A _03576_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_687 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07091_ _00355_ VGND VGND VPWR VPWR _00366_ sky130_fd_sc_hd__buf_4
XANTENNA__12392__A _01517_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11898__A1 _06428_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11898__B2 _06439_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09801_ _01782_ _01784_ _01990_ VGND VGND VPWR VPWR _01991_ sky130_fd_sc_hd__o21a_1
XFILLER_0_10_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07993_ _00035_ _00036_ VGND VGND VPWR VPWR _00037_ sky130_fd_sc_hd__nand2_1
X_09732_ _01541_ _01543_ _01692_ _01914_ VGND VGND VPWR VPWR _01915_ sky130_fd_sc_hd__a31o_2
XANTENNA__12311__A2 _00575_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09663_ _00670_ _00145_ VGND VGND VPWR VPWR _01839_ sky130_fd_sc_hd__nand2_1
XANTENNA__11455__B _02673_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07652__C _06472_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08614_ _00500_ _00502_ _00691_ VGND VGND VPWR VPWR _00692_ sky130_fd_sc_hd__o21a_1
XANTENNA__08467__D _05203_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09594_ _03510_ _03762_ VGND VGND VPWR VPWR _01764_ sky130_fd_sc_hd__nand2_1
XTAP_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08545_ _00614_ _00615_ VGND VGND VPWR VPWR _00616_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08476_ _00340_ _00540_ VGND VGND VPWR VPWR _00542_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_77_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07427_ net40 VGND VGND VPWR VPWR _04048_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_147_486 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13024__B1 _05515_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_648 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07358_ _01295_ _02664_ _02719_ _01306_ VGND VGND VPWR VPWR _03290_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07289_ net62 net12 net61 _00869_ VGND VGND VPWR VPWR _02532_ sky130_fd_sc_hd__and4_1
XANTENNA__10815__A _06937_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09028_ _00998_ _01002_ _01143_ VGND VGND VPWR VPWR _01145_ sky130_fd_sc_hd__nand3_1
XANTENNA__07396__A _03696_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11349__C _01956_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11646__A _02249_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12838__B1 _02727_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14022__A _05424_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13990_ _06558_ _06575_ VGND VGND VPWR VPWR _06576_ sky130_fd_sc_hd__xnor2_1
X_12941_ _04570_ _04571_ _02699_ VGND VGND VPWR VPWR _05440_ sky130_fd_sc_hd__a21o_1
XTAP_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12872_ _05239_ _05240_ VGND VGND VPWR VPWR _05364_ sky130_fd_sc_hd__or2b_1
XTAP_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11823_ _04208_ _04209_ VGND VGND VPWR VPWR _04210_ sky130_fd_sc_hd__nor2_1
XANTENNA__13580__B _03783_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12477__A _04714_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10616__A2 _01060_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11754_ _04124_ _04133_ VGND VGND VPWR VPWR _04134_ sky130_fd_sc_hd__xor2_1
XTAP_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10705_ _02968_ _02969_ VGND VGND VPWR VPWR _02981_ sky130_fd_sc_hd__or2_1
XTAP_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11685_ _04055_ _02608_ _04056_ VGND VGND VPWR VPWR _04058_ sky130_fd_sc_hd__a21o_1
XFILLER_0_102_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13424_ _05413_ _05852_ _05953_ VGND VGND VPWR VPWR _05954_ sky130_fd_sc_hd__and3_1
X_10636_ _02865_ _02892_ VGND VGND VPWR VPWR _02906_ sky130_fd_sc_hd__nor2_1
XANTENNA__09234__A2 _01368_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13355_ _05875_ _05877_ VGND VGND VPWR VPWR _05878_ sky130_fd_sc_hd__or2_1
XFILLER_0_140_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10567_ _02826_ _02829_ VGND VGND VPWR VPWR _02830_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_140_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13824__A1_N _03414_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12306_ _01400_ _01780_ VGND VGND VPWR VPWR _04742_ sky130_fd_sc_hd__nand2_1
X_13286_ _05788_ _05807_ VGND VGND VPWR VPWR _05809_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10498_ _02749_ _02753_ VGND VGND VPWR VPWR _02754_ sky130_fd_sc_hd__and2b_1
X_12237_ _04651_ _04650_ VGND VGND VPWR VPWR _04666_ sky130_fd_sc_hd__and2b_1
X_12168_ _04519_ _04530_ VGND VGND VPWR VPWR _04590_ sky130_fd_sc_hd__nor2_1
XANTENNA__11556__A _00497_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11119_ _03429_ _03421_ VGND VGND VPWR VPWR _03437_ sky130_fd_sc_hd__and2b_1
X_12099_ _04511_ _04513_ VGND VGND VPWR VPWR _04514_ sky130_fd_sc_hd__xor2_2
Xinput6 a[14] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__buf_4
XFILLER_0_36_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08330_ _00464_ _00376_ _00381_ _02051_ VGND VGND VPWR VPWR _00382_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_52_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_475 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08261_ _00304_ _00305_ _02018_ _00143_ VGND VGND VPWR VPWR _00306_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_6_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07212_ _01525_ _01492_ VGND VGND VPWR VPWR _01689_ sky130_fd_sc_hd__xor2_1
XFILLER_0_144_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08192_ _00194_ _00235_ VGND VGND VPWR VPWR _00236_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07143_ net1 _00923_ net61 net60 VGND VGND VPWR VPWR _00934_ sky130_fd_sc_hd__and4_1
XFILLER_0_6_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12780__A2 _02849_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10791__A1 _02149_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10791__B2 _02105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08736__A1 _00377_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08736__B2 _02993_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07976_ _07021_ _07026_ VGND VGND VPWR VPWR _00020_ sky130_fd_sc_hd__nand2_1
X_09715_ _06483_ _00607_ _01892_ _01894_ VGND VGND VPWR VPWR _01896_ sky130_fd_sc_hd__and4_1
XANTENNA__11099__A2 _01066_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12296__A1 _02427_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12296__B2 _02188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09161__A1 _03070_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09161__B2 _02456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09646_ _01807_ _01820_ VGND VGND VPWR VPWR _01822_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_96_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11913__B _00159_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09577_ _01738_ _01742_ VGND VGND VPWR VPWR _01746_ sky130_fd_sc_hd__nor2_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08528_ _00596_ _00597_ VGND VGND VPWR VPWR _00598_ sky130_fd_sc_hd__and2_2
XANTENNA__12599__A2 _01059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08459_ _00496_ _00522_ VGND VGND VPWR VPWR _00523_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_53_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11470_ _03819_ _03821_ VGND VGND VPWR VPWR _03822_ sky130_fd_sc_hd__and2b_1
XFILLER_0_18_484 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12744__B _03681_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10421_ _02127_ _02459_ VGND VGND VPWR VPWR _02670_ sky130_fd_sc_hd__nand2_1
XANTENNA__07838__B _01350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08975__A1 _05577_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13140_ _05652_ _05653_ _05658_ VGND VGND VPWR VPWR _05659_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_103_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10352_ _02433_ VGND VGND VPWR VPWR _02594_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10782__A1 _06637_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10782__B2 _06937_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13071_ _02483_ _02484_ _02485_ _02486_ VGND VGND VPWR VPWR _05583_ sky130_fd_sc_hd__a211o_1
X_10283_ _02318_ _02516_ VGND VGND VPWR VPWR _02518_ sky130_fd_sc_hd__or2_1
X_12022_ _06626_ _06450_ _03683_ _03679_ VGND VGND VPWR VPWR _04429_ sky130_fd_sc_hd__and4_1
XANTENNA__08669__B net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09491__D net52 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13973_ _06157_ _06159_ VGND VGND VPWR VPWR _06557_ sky130_fd_sc_hd__or2_1
X_12924_ _04629_ _05316_ _05420_ VGND VGND VPWR VPWR _05421_ sky130_fd_sc_hd__o21a_1
XANTENNA__07933__A1_N _01470_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12855_ _01584_ _01412_ VGND VGND VPWR VPWR _05345_ sky130_fd_sc_hd__nand2_1
XTAP_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_716 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11806_ _04185_ _04190_ VGND VGND VPWR VPWR _04192_ sky130_fd_sc_hd__xor2_1
XTAP_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12786_ _01585_ _01059_ VGND VGND VPWR VPWR _05270_ sky130_fd_sc_hd__nand2_1
XTAP_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_855 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11737_ _04083_ _04115_ VGND VGND VPWR VPWR _04116_ sky130_fd_sc_hd__and2_1
XFILLER_0_138_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12217__A2_N _03750_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11668_ _04038_ _04039_ VGND VGND VPWR VPWR _04040_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_126_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13407_ _05932_ _05935_ VGND VGND VPWR VPWR _05936_ sky130_fd_sc_hd__and2_1
XFILLER_0_52_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10619_ _02885_ _02886_ VGND VGND VPWR VPWR _02887_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07748__B _06873_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11599_ _03961_ _03963_ VGND VGND VPWR VPWR _03964_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13338_ _05855_ _05859_ VGND VGND VPWR VPWR _05860_ sky130_fd_sc_hd__xor2_1
XFILLER_0_110_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13269_ _05787_ _05778_ VGND VGND VPWR VPWR _05793_ sky130_fd_sc_hd__nor2_1
XFILLER_0_121_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07830_ _06957_ _06958_ VGND VGND VPWR VPWR _06959_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07483__B _04367_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07761_ _06884_ _06888_ _06889_ VGND VGND VPWR VPWR _06890_ sky130_fd_sc_hd__a21bo_1
X_09500_ _01552_ _01660_ VGND VGND VPWR VPWR _01661_ sky130_fd_sc_hd__and2_1
X_07692_ _06820_ VGND VGND VPWR VPWR _06821_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09431_ _01272_ VGND VGND VPWR VPWR _01586_ sky130_fd_sc_hd__buf_4
XFILLER_0_78_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_340 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09362_ _01350_ _01505_ _01509_ VGND VGND VPWR VPWR _01510_ sky130_fd_sc_hd__and3_1
XFILLER_0_75_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08313_ _00202_ _00203_ _06998_ VGND VGND VPWR VPWR _00363_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_129_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09293_ _00899_ _01053_ VGND VGND VPWR VPWR _01435_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08244_ _00132_ _00133_ VGND VGND VPWR VPWR _00288_ sky130_fd_sc_hd__and2b_1
XFILLER_0_145_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08175_ _06845_ _00218_ VGND VGND VPWR VPWR _00219_ sky130_fd_sc_hd__or2_2
XFILLER_0_6_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07126_ _00737_ _00726_ VGND VGND VPWR VPWR _00748_ sky130_fd_sc_hd__and2b_1
XFILLER_0_113_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12580__A _03740_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07674__A net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07959_ _06765_ VGND VGND VPWR VPWR _00003_ sky130_fd_sc_hd__clkbuf_4
X_10970_ _04862_ _00604_ _01506_ _04873_ VGND VGND VPWR VPWR _03273_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09629_ _01801_ _01802_ VGND VGND VPWR VPWR _01803_ sky130_fd_sc_hd__and2b_1
XFILLER_0_85_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12640_ _00915_ _02855_ VGND VGND VPWR VPWR _05109_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_310 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12571_ _04991_ _04993_ _05031_ _05032_ VGND VGND VPWR VPWR _05033_ sky130_fd_sc_hd__a31o_1
XFILLER_0_81_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11522_ _03826_ _03832_ VGND VGND VPWR VPWR _03879_ sky130_fd_sc_hd__xor2_1
XFILLER_0_19_771 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07999__A2 _04917_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12992__A2 _05494_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07568__B _05588_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11453_ _03801_ _03802_ _03532_ _03681_ VGND VGND VPWR VPWR _03803_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_80_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_251 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10404_ _02007_ _02117_ VGND VGND VPWR VPWR _02651_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14172_ _06616_ _06642_ _06753_ _05841_ VGND VGND VPWR VPWR _06772_ sky130_fd_sc_hd__or4b_4
X_11384_ _03725_ _03726_ VGND VGND VPWR VPWR _03727_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10755__A1 _00526_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13123_ _05215_ _05171_ _05212_ VGND VGND VPWR VPWR _05640_ sky130_fd_sc_hd__or3_1
XFILLER_0_0_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10335_ _02372_ _02573_ VGND VGND VPWR VPWR _02575_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13054_ _05551_ _05554_ VGND VGND VPWR VPWR _05564_ sky130_fd_sc_hd__and2_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10266_ _02342_ VGND VGND VPWR VPWR _02500_ sky130_fd_sc_hd__inv_2
XANTENNA__11818__B _03682_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12005_ _00843_ _02090_ _02088_ _00844_ VGND VGND VPWR VPWR _04410_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_84_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10197_ _02087_ _02097_ VGND VGND VPWR VPWR _02425_ sky130_fd_sc_hd__and2b_1
X_13956_ _06477_ _06465_ VGND VGND VPWR VPWR _06539_ sky130_fd_sc_hd__and2b_1
XFILLER_0_88_424 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12649__B _01061_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12907_ _05399_ _05402_ VGND VGND VPWR VPWR _05403_ sky130_fd_sc_hd__xor2_1
X_13887_ _06462_ _06448_ _06447_ VGND VGND VPWR VPWR _06463_ sky130_fd_sc_hd__o21a_1
XFILLER_0_75_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10145__A1_N _05027_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08565__D _04939_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12838_ _00742_ _02724_ _02727_ _00392_ VGND VGND VPWR VPWR _05327_ sky130_fd_sc_hd__a22oi_2
XTAP_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10169__B _00741_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11235__A2 _01062_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12769_ _05232_ _05250_ VGND VGND VPWR VPWR _05251_ sky130_fd_sc_hd__xor2_1
XFILLER_0_29_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07759__A _00453_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08581__C _06765_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput20 a[27] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_4
Xinput31 a[8] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__buf_2
XFILLER_0_142_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput42 b[18] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_448 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput53 b[28] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_4_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput64 b[9] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__buf_4
XFILLER_0_12_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12735__A2 _05150_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09980_ _01664_ VGND VGND VPWR VPWR _02187_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_110_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08931_ _01037_ _00870_ _01038_ VGND VGND VPWR VPWR _01039_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_110_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08862_ _00961_ _00962_ VGND VGND VPWR VPWR _00963_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08102__B _00145_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07813_ _06940_ _06941_ VGND VGND VPWR VPWR _06942_ sky130_fd_sc_hd__and2b_1
X_08793_ _00886_ _00887_ VGND VGND VPWR VPWR _00888_ sky130_fd_sc_hd__and2b_1
XANTENNA__13448__B1 _02731_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07744_ _06819_ VGND VGND VPWR VPWR _06873_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08756__C _00846_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07678__A1 _00442_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07675_ _00442_ _00989_ _06733_ _06744_ VGND VGND VPWR VPWR _06755_ sky130_fd_sc_hd__and4_1
XANTENNA__07678__B2 _02051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09414_ _04510_ _00661_ net17 net18 VGND VGND VPWR VPWR _01567_ sky130_fd_sc_hd__and4_1
XANTENNA__10079__B _02293_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_855 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09345_ _01409_ _01420_ _01365_ VGND VGND VPWR VPWR _01491_ sky130_fd_sc_hd__a21o_1
XFILLER_0_90_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09276_ _02051_ _01062_ _01415_ _00464_ VGND VGND VPWR VPWR _01417_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_63_847 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08227_ _00269_ _00270_ VGND VGND VPWR VPWR _00271_ sky130_fd_sc_hd__and2b_1
XANTENNA__07388__B _03609_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10095__A net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08158_ _00190_ _00191_ _00201_ VGND VGND VPWR VPWR _00202_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_43_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07109_ net27 VGND VGND VPWR VPWR _00563_ sky130_fd_sc_hd__buf_6
X_08089_ _00007_ _00036_ _00035_ VGND VGND VPWR VPWR _00133_ sky130_fd_sc_hd__a21bo_1
XANTENNA__12741__C _02133_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10120_ _02336_ _02201_ _02339_ VGND VGND VPWR VPWR _02340_ sky130_fd_sc_hd__nor3_1
X_10051_ _02263_ _02264_ VGND VGND VPWR VPWR _02265_ sky130_fd_sc_hd__nand2_1
XANTENNA__09108__B _01232_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13853__B _03679_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13810_ _02189_ _01955_ _03686_ _02188_ VGND VGND VPWR VPWR _06378_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_97_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13741_ _02090_ _02855_ VGND VGND VPWR VPWR _06302_ sky130_fd_sc_hd__nand2_1
XANTENNA__09124__A _01248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10953_ _00298_ _00608_ VGND VGND VPWR VPWR _03254_ sky130_fd_sc_hd__nand2_1
XANTENNA__08330__A2 _00376_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13672_ _06221_ _06224_ _06225_ VGND VGND VPWR VPWR _06226_ sky130_fd_sc_hd__a21o_1
XFILLER_0_39_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10884_ _03137_ _03177_ VGND VGND VPWR VPWR _03178_ sky130_fd_sc_hd__nor2_1
XANTENNA__08963__A _04169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12623_ _05085_ _05088_ _05089_ VGND VGND VPWR VPWR _05090_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_109_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12485__A _00784_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09778__B net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12554_ _05010_ _05012_ _05013_ VGND VGND VPWR VPWR _05014_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_53_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11505_ _03858_ _03853_ _03857_ VGND VGND VPWR VPWR _03860_ sky130_fd_sc_hd__and3_1
XFILLER_0_123_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12485_ _00784_ _00779_ _00742_ _00741_ VGND VGND VPWR VPWR _04938_ sky130_fd_sc_hd__nand4_1
XFILLER_0_108_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14224_ _00406_ _00408_ VGND VGND VPWR VPWR _06808_ sky130_fd_sc_hd__nor2_1
X_11436_ _03750_ VGND VGND VPWR VPWR _03785_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_123_256 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12932__B _05429_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14155_ _05960_ _06753_ VGND VGND VPWR VPWR _06754_ sky130_fd_sc_hd__nor2_1
XANTENNA__13390__A2 _03681_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11367_ _03693_ _03695_ _03706_ VGND VGND VPWR VPWR _03709_ sky130_fd_sc_hd__nor3_1
X_13106_ _05608_ _05620_ VGND VGND VPWR VPWR _05622_ sky130_fd_sc_hd__and2_1
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10318_ _02552_ _02556_ VGND VGND VPWR VPWR _02557_ sky130_fd_sc_hd__xor2_1
X_14086_ _06678_ _06679_ VGND VGND VPWR VPWR _06681_ sky130_fd_sc_hd__nor2_2
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11298_ _02910_ _03630_ _03633_ VGND VGND VPWR VPWR _03634_ sky130_fd_sc_hd__o21a_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13037_ _05543_ _05545_ VGND VGND VPWR VPWR _05546_ sky130_fd_sc_hd__and2b_2
X_10249_ _02480_ _02481_ VGND VGND VPWR VPWR _02482_ sky130_fd_sc_hd__or2_4
XFILLER_0_119_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_700 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08857__B _04169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13939_ _06518_ _06519_ VGND VGND VPWR VPWR _06520_ sky130_fd_sc_hd__and2b_1
XFILLER_0_44_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07460_ _01470_ _04378_ _04389_ net164 VGND VGND VPWR VPWR _04411_ sky130_fd_sc_hd__a31o_1
XFILLER_0_29_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07391_ _02949_ _03631_ VGND VGND VPWR VPWR _03653_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12395__A _00782_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09130_ _01253_ _01255_ VGND VGND VPWR VPWR _01256_ sky130_fd_sc_hd__and2_1
XFILLER_0_60_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09061_ _01180_ VGND VGND VPWR VPWR _01181_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_60_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08012_ _06921_ _07053_ _07052_ VGND VGND VPWR VPWR _00056_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_13_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_73 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09963_ net54 VGND VGND VPWR VPWR _02168_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__08113__A _01361_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08914_ _01018_ _01019_ VGND VGND VPWR VPWR _01020_ sky130_fd_sc_hd__nand2_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09894_ _06626_ _06450_ _02090_ _02088_ VGND VGND VPWR VPWR _02092_ sky130_fd_sc_hd__and4_1
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08845_ _00563_ _00639_ _04180_ _04191_ VGND VGND VPWR VPWR _00944_ sky130_fd_sc_hd__and4_1
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08767__B _00859_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08776_ _00496_ _00522_ _00867_ _00868_ VGND VGND VPWR VPWR _00870_ sky130_fd_sc_hd__a31oi_4
X_07727_ _06851_ _06854_ _06855_ VGND VGND VPWR VPWR _06856_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_95_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07658_ _05934_ _06318_ _06296_ VGND VGND VPWR VPWR _06571_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_67_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07589_ _05445_ _05467_ _02105_ _00650_ VGND VGND VPWR VPWR _05818_ sky130_fd_sc_hd__and4_1
XFILLER_0_137_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09328_ _01472_ VGND VGND VPWR VPWR _01473_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10537__B _00293_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09259_ _01396_ _01397_ VGND VGND VPWR VPWR _01398_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_543 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12270_ _03414_ _01181_ _01250_ _01066_ VGND VGND VPWR VPWR _04702_ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11221_ _03545_ _03547_ _03546_ VGND VGND VPWR VPWR _03549_ sky130_fd_sc_hd__nand3_2
XANTENNA__10553__A _00377_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_790 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11383__A1 _02246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11383__B2 _02249_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11152_ _03245_ _03472_ VGND VGND VPWR VPWR _03473_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_462 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10103_ _02311_ _02320_ VGND VGND VPWR VPWR _02321_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10703__D _01412_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11083_ _03276_ _03277_ VGND VGND VPWR VPWR _03397_ sky130_fd_sc_hd__or2_1
XANTENNA__07339__B1 _02171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10034_ _00843_ VGND VGND VPWR VPWR _02246_ sky130_fd_sc_hd__buf_4
X_11985_ _04357_ _04385_ _04386_ _04387_ VGND VGND VPWR VPWR _04388_ sky130_fd_sc_hd__nand4_1
XANTENNA_output118_A net118 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10936_ _03230_ _03229_ VGND VGND VPWR VPWR _03236_ sky130_fd_sc_hd__or2_1
X_13724_ _06281_ _06282_ VGND VGND VPWR VPWR _06283_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13655_ _05976_ VGND VGND VPWR VPWR _06207_ sky130_fd_sc_hd__inv_2
X_10867_ _03156_ _03157_ VGND VGND VPWR VPWR _03160_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12606_ _05051_ _05047_ VGND VGND VPWR VPWR _05072_ sky130_fd_sc_hd__xor2_1
XFILLER_0_94_791 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13586_ _06018_ _05985_ _06121_ _06129_ VGND VGND VPWR VPWR _06132_ sky130_fd_sc_hd__a31o_1
XFILLER_0_27_847 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10798_ _06461_ _02168_ VGND VGND VPWR VPWR _03084_ sky130_fd_sc_hd__nand2_1
XPHY_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07102__A _00475_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12537_ _04986_ _04995_ VGND VGND VPWR VPWR _04996_ sky130_fd_sc_hd__xor2_1
XFILLER_0_53_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12468_ _04900_ _04902_ VGND VGND VPWR VPWR _04920_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09955__C _02158_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14207_ _01766_ _01777_ VGND VGND VPWR VPWR _06798_ sky130_fd_sc_hd__and2_1
XANTENNA__11559__A _00486_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11419_ _06775_ _03744_ VGND VGND VPWR VPWR _03766_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12399_ _04842_ _04843_ VGND VGND VPWR VPWR _04844_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_22_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14138_ _06708_ _06735_ VGND VGND VPWR VPWR _06736_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14069_ _06078_ _02743_ _02742_ _06075_ VGND VGND VPWR VPWR _06662_ sky130_fd_sc_hd__a22oi_1
XANTENNA__09971__B _02149_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11677__A2 _03773_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08630_ _00707_ _00709_ VGND VGND VPWR VPWR _00710_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_146_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08561_ _00527_ _00632_ _00633_ VGND VGND VPWR VPWR _00634_ sky130_fd_sc_hd__a21o_1
XANTENNA__12626__A1 _01413_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07512_ _04840_ _04961_ _04972_ VGND VGND VPWR VPWR _04983_ sky130_fd_sc_hd__o21bai_2
X_08492_ _00463_ _00558_ VGND VGND VPWR VPWR _00559_ sky130_fd_sc_hd__nor2_2
XFILLER_0_49_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07443_ _04202_ _04213_ VGND VGND VPWR VPWR _04224_ sky130_fd_sc_hd__and2b_1
XFILLER_0_119_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10638__A _00859_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07374_ _02839_ _03444_ _03433_ VGND VGND VPWR VPWR _03466_ sky130_fd_sc_hd__o21a_1
XFILLER_0_18_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08108__A _05478_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10357__B _00101_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09113_ _01234_ _01237_ VGND VGND VPWR VPWR _01238_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_45_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12853__A _00572_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09044_ _01113_ _01114_ _01161_ VGND VGND VPWR VPWR _01162_ sky130_fd_sc_hd__a21o_1
XFILLER_0_72_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09865__C _03707_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09558__A1 _00844_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_861 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09558__B2 _00843_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10092__B _02308_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09881__B _00486_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09946_ _02056_ _02037_ _02038_ _02148_ VGND VGND VPWR VPWR _02150_ sky130_fd_sc_hd__o31ai_4
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09877_ _02059_ _02060_ _02073_ VGND VGND VPWR VPWR _02074_ sky130_fd_sc_hd__a21o_1
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08828_ _00901_ net11 VGND VGND VPWR VPWR _00926_ sky130_fd_sc_hd__and2_1
XTAP_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08759_ _00676_ _00681_ _00850_ VGND VGND VPWR VPWR _00851_ sky130_fd_sc_hd__nor3_1
XFILLER_0_68_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11932__A _00114_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11770_ _05445_ _05731_ _01246_ net19 VGND VGND VPWR VPWR _04152_ sky130_fd_sc_hd__and4_1
XTAP_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12747__B _03678_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10721_ _02997_ _02990_ _02995_ VGND VGND VPWR VPWR _02999_ sky130_fd_sc_hd__and3_1
XTAP_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13440_ _05970_ VGND VGND VPWR VPWR _05971_ sky130_fd_sc_hd__inv_2
X_10652_ _02922_ _02890_ VGND VGND VPWR VPWR _02923_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09246__B1 _00613_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09797__A1 _03070_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_510 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13371_ _05360_ _05895_ VGND VGND VPWR VPWR _05896_ sky130_fd_sc_hd__nand2_1
X_10583_ _02845_ _02846_ VGND VGND VPWR VPWR _02847_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12322_ _04750_ _04756_ _04758_ VGND VGND VPWR VPWR _04759_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_106_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07272__A2 _02335_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12253_ _04677_ _04682_ VGND VGND VPWR VPWR _04683_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_50_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11204_ net178 _03528_ _03529_ VGND VGND VPWR VPWR _03530_ sky130_fd_sc_hd__nor3_1
X_12184_ _03608_ _03578_ _03610_ VGND VGND VPWR VPWR _04607_ sky130_fd_sc_hd__or3b_1
XFILLER_0_102_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11135_ _03002_ _03453_ VGND VGND VPWR VPWR _03454_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07592__A _02007_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11066_ _03375_ _03377_ VGND VGND VPWR VPWR _03379_ sky130_fd_sc_hd__nand2_1
X_10017_ _02222_ _02227_ VGND VGND VPWR VPWR _02228_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08288__A1 _00497_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11968_ _04296_ net144 _04368_ VGND VGND VPWR VPWR _04370_ sky130_fd_sc_hd__nor3_1
XFILLER_0_25_89 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13707_ _02726_ _05887_ _06264_ VGND VGND VPWR VPWR _06265_ sky130_fd_sc_hd__a21bo_1
X_10919_ _02171_ _02758_ _02720_ _02467_ VGND VGND VPWR VPWR _03217_ sky130_fd_sc_hd__a22oi_1
X_11899_ _04292_ _04293_ _03059_ _03682_ VGND VGND VPWR VPWR _04294_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_129_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13638_ _06188_ VGND VGND VPWR VPWR _06189_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10177__B _06733_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_761 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09966__B _00989_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_143_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13569_ _06102_ _06111_ _06112_ VGND VGND VPWR VPWR _06113_ sky130_fd_sc_hd__o21a_1
XFILLER_0_125_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_699 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12792__B1 _02727_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07090_ net31 VGND VGND VPWR VPWR _00355_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_140_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12392__B _01780_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09982__A _01505_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11898__A2 _01954_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09800_ _01982_ _01989_ VGND VGND VPWR VPWR _01990_ sky130_fd_sc_hd__xnor2_1
X_07992_ _07030_ _00034_ VGND VGND VPWR VPWR _00036_ sky130_fd_sc_hd__or2_1
XFILLER_0_66_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09731_ _01539_ _01693_ _01913_ _01691_ VGND VGND VPWR VPWR _01914_ sky130_fd_sc_hd__a31o_1
X_09662_ _01740_ _01741_ VGND VGND VPWR VPWR _01838_ sky130_fd_sc_hd__nor2_1
XANTENNA__07652__D _06494_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08371__A1_N _01744_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08613_ _00689_ _00690_ VGND VGND VPWR VPWR _00691_ sky130_fd_sc_hd__nor2_1
X_09593_ _03685_ _01761_ _01762_ VGND VGND VPWR VPWR _01763_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_77_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08544_ _01372_ _04268_ _00612_ _00613_ VGND VGND VPWR VPWR _00615_ sky130_fd_sc_hd__nand4_1
XTAP_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08475_ _00538_ _00539_ VGND VGND VPWR VPWR _00540_ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07426_ _04026_ VGND VGND VPWR VPWR _04037_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_58_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13024__B2 _05513_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07357_ _01744_ _03268_ _02697_ _02686_ VGND VGND VPWR VPWR _03279_ sky130_fd_sc_hd__a31o_1
XFILLER_0_134_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12583__A _00745_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_90 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07677__A _06744_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07288_ _00891_ _01000_ _01055_ _01033_ VGND VGND VPWR VPWR _02521_ sky130_fd_sc_hd__a31o_1
XANTENNA__10815__B _02735_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_142_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09027_ _00998_ _01002_ _01143_ VGND VGND VPWR VPWR _01144_ sky130_fd_sc_hd__a21o_1
XFILLER_0_13_360 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09892__A _01601_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09951__A1 _01339_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12838__A1 _00742_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09929_ _02129_ _02112_ _02113_ VGND VGND VPWR VPWR _02131_ sky130_fd_sc_hd__nand3_1
XANTENNA__08301__A _04004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12838__B2 _00392_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12940_ _04573_ _05437_ _05438_ VGND VGND VPWR VPWR _05439_ sky130_fd_sc_hd__a21o_1
XFILLER_0_99_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12871_ _05255_ _05257_ _05254_ VGND VGND VPWR VPWR _05363_ sky130_fd_sc_hd__a21oi_1
XTAP_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11662__A _00258_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11822_ _04207_ _04203_ _04204_ VGND VGND VPWR VPWR _04209_ sky130_fd_sc_hd__nor3_1
XTAP_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12477__B _02008_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11753_ _04127_ _04131_ _04132_ VGND VGND VPWR VPWR _04133_ sky130_fd_sc_hd__o21bai_1
XTAP_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10704_ _02978_ _02979_ VGND VGND VPWR VPWR _02980_ sky130_fd_sc_hd__nand2_1
XTAP_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11684_ _04055_ _02608_ _04056_ VGND VGND VPWR VPWR _04057_ sky130_fd_sc_hd__and3_1
XTAP_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__14212__B1 _00344_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10635_ _02853_ _02864_ VGND VGND VPWR VPWR _02904_ sky130_fd_sc_hd__and2b_1
XFILLER_0_102_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13423_ _05948_ _05952_ VGND VGND VPWR VPWR _05953_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_107_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13354_ _05876_ _05874_ VGND VGND VPWR VPWR _05877_ sky130_fd_sc_hd__nor2_1
X_10566_ _02805_ _02827_ VGND VGND VPWR VPWR _02829_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12305_ _04727_ _04726_ VGND VGND VPWR VPWR _04740_ sky130_fd_sc_hd__and2b_1
X_13285_ _05472_ _05491_ _05725_ _05732_ VGND VGND VPWR VPWR _05807_ sky130_fd_sc_hd__and4_2
X_10497_ _01473_ _02721_ _02750_ _02752_ VGND VGND VPWR VPWR _02753_ sky130_fd_sc_hd__a31o_1
X_12236_ _00375_ _03750_ _04662_ _04663_ VGND VGND VPWR VPWR _04665_ sky130_fd_sc_hd__a31o_1
X_12167_ _04534_ _04535_ VGND VGND VPWR VPWR _04589_ sky130_fd_sc_hd__and2_1
X_11118_ _03423_ _03435_ VGND VGND VPWR VPWR _03436_ sky130_fd_sc_hd__xnor2_2
XANTENNA__11556__B _02120_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12098_ _04382_ _04383_ _04384_ _04442_ _04512_ VGND VGND VPWR VPWR _04513_ sky130_fd_sc_hd__a41o_2
X_11049_ _03351_ _03359_ VGND VGND VPWR VPWR _03360_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput7 a[15] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_4
XFILLER_0_36_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08260_ _00138_ _04906_ _04928_ _06417_ VGND VGND VPWR VPWR _00305_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_117_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_430 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_487 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07211_ _01656_ _01667_ VGND VGND VPWR VPWR _01678_ sky130_fd_sc_hd__nand2_1
XFILLER_0_116_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08191_ _00196_ _00198_ VGND VGND VPWR VPWR _00235_ sky130_fd_sc_hd__xor2_1
XFILLER_0_144_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_794 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07142_ net12 VGND VGND VPWR VPWR _00923_ sky130_fd_sc_hd__buf_6
XFILLER_0_15_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10791__A2 net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08736__A2 _00114_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07975_ _00016_ _00018_ VGND VGND VPWR VPWR _00019_ sky130_fd_sc_hd__xor2_1
X_09714_ _06494_ _00608_ _01892_ _01894_ VGND VGND VPWR VPWR _01895_ sky130_fd_sc_hd__a22oi_1
XANTENNA__12296__A2 _02190_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07960__A _00003_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09161__A2 _01188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09645_ _01818_ _01819_ VGND VGND VPWR VPWR _01820_ sky130_fd_sc_hd__or2_2
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09576_ _01743_ VGND VGND VPWR VPWR _01745_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11913__C _03683_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08527_ _00570_ _00594_ VGND VGND VPWR VPWR _00597_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10098__A _04081_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08458_ _00520_ _00521_ VGND VGND VPWR VPWR _00522_ sky130_fd_sc_hd__nor2_2
XFILLER_0_65_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07409_ _01197_ VGND VGND VPWR VPWR _03850_ sky130_fd_sc_hd__buf_2
XFILLER_0_18_463 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08389_ _00880_ _04180_ _04191_ _04169_ VGND VGND VPWR VPWR _00446_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10420_ net21 _02667_ _02668_ VGND VGND VPWR VPWR _02669_ sky130_fd_sc_hd__a21bo_1
XANTENNA__07838__C _06965_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08975__A2 _00373_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10351_ _02496_ _02498_ _02591_ VGND VGND VPWR VPWR _02593_ sky130_fd_sc_hd__nand3_1
XFILLER_0_21_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10782__A2 _02726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13070_ _02491_ _02713_ VGND VGND VPWR VPWR _05582_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10282_ _02318_ _02516_ VGND VGND VPWR VPWR _02517_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12021_ _04369_ _04371_ VGND VGND VPWR VPWR _04428_ sky130_fd_sc_hd__and2b_1
XANTENNA__08669__C net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08388__D net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13972_ _06553_ _06555_ VGND VGND VPWR VPWR _06556_ sky130_fd_sc_hd__nor2_1
XANTENNA__08966__A _04268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12923_ _05318_ _05419_ VGND VGND VPWR VPWR _05420_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12488__A _01518_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11392__A _00112_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12854_ _05342_ _05343_ VGND VGND VPWR VPWR _05344_ sky130_fd_sc_hd__nor2_1
XTAP_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11805_ _02466_ _02679_ _04188_ _04189_ VGND VGND VPWR VPWR _04190_ sky130_fd_sc_hd__o31a_1
XFILLER_0_139_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_739 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12785_ _01586_ _01059_ _05092_ _05267_ VGND VGND VPWR VPWR _05268_ sky130_fd_sc_hd__a31o_1
XFILLER_0_95_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11736_ _04061_ _04082_ VGND VGND VPWR VPWR _04115_ sky130_fd_sc_hd__or2_1
XTAP_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11667_ _00004_ _06885_ _00416_ _01288_ VGND VGND VPWR VPWR _04039_ sky130_fd_sc_hd__and4_1
X_13406_ _05933_ VGND VGND VPWR VPWR _05935_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10618_ _00635_ _04939_ _01060_ _01413_ VGND VGND VPWR VPWR _02886_ sky130_fd_sc_hd__and4_1
XFILLER_0_113_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11598_ _03941_ _03962_ VGND VGND VPWR VPWR _03963_ sky130_fd_sc_hd__or2_1
XFILLER_0_107_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07110__A net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10549_ _02807_ _02808_ _02809_ VGND VGND VPWR VPWR _02810_ sky130_fd_sc_hd__and3_1
X_13337_ _05856_ _05858_ VGND VGND VPWR VPWR _05859_ sky130_fd_sc_hd__nand2_1
XFILLER_0_106_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13268_ _05787_ _05792_ VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__xnor2_4
XANTENNA__09915__A1 _02138_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11567__A _03532_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12219_ _00459_ _00608_ _01180_ _01249_ VGND VGND VPWR VPWR _04646_ sky130_fd_sc_hd__nand4_4
XFILLER_0_110_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10471__A _02723_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13199_ _05719_ _05722_ _05723_ VGND VGND VPWR VPWR _05724_ sky130_fd_sc_hd__a21oi_2
XANTENNA__09037__A _00544_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07760_ _00442_ _06775_ _06887_ VGND VGND VPWR VPWR _06889_ sky130_fd_sc_hd__a21o_1
XANTENNA__10289__A1 _05742_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10289__B2 _00628_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07691_ net34 VGND VGND VPWR VPWR _06820_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__07154__A1 net1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12398__A _00374_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07154__B2 net61 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09430_ _01584_ VGND VGND VPWR VPWR _01585_ sky130_fd_sc_hd__buf_4
XFILLER_0_59_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09361_ _01383_ _01508_ VGND VGND VPWR VPWR _01509_ sky130_fd_sc_hd__nand2_1
X_08312_ _00204_ _00205_ _00361_ VGND VGND VPWR VPWR _00362_ sky130_fd_sc_hd__or3_4
XFILLER_0_86_171 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09292_ _01054_ _01239_ VGND VGND VPWR VPWR _01434_ sky130_fd_sc_hd__or2_4
XFILLER_0_129_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08243_ _00285_ _00286_ VGND VGND VPWR VPWR _00287_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_411 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08174_ _03598_ _06844_ VGND VGND VPWR VPWR _00218_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09603__B1 _00574_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08116__A _00159_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07125_ net27 _00705_ net28 _00573_ VGND VGND VPWR VPWR _00737_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_61 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_447 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07955__A _03532_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12580__B _00742_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07917__B1 _04367_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07958_ _00000_ _00001_ VGND VGND VPWR VPWR _00002_ sky130_fd_sc_hd__and2_1
XANTENNA__07690__A _06818_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_403 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07889_ _06961_ _07017_ VGND VGND VPWR VPWR _07018_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09628_ _01800_ _01796_ VGND VGND VPWR VPWR _01802_ sky130_fd_sc_hd__or2b_1
X_09559_ _01724_ _01725_ _00654_ _01472_ VGND VGND VPWR VPWR _01726_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_65_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12570_ _04929_ _04990_ VGND VGND VPWR VPWR _05032_ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11521_ _03772_ _03778_ VGND VGND VPWR VPWR _03878_ sky130_fd_sc_hd__xor2_1
XFILLER_0_136_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11452_ _06964_ _01953_ _02134_ _06966_ VGND VGND VPWR VPWR _03802_ sky130_fd_sc_hd__a22oi_1
X_10403_ _01178_ _02648_ _02649_ VGND VGND VPWR VPWR _02650_ sky130_fd_sc_hd__a21bo_1
X_14171_ _06750_ _06770_ VGND VGND VPWR VPWR _06771_ sky130_fd_sc_hd__xnor2_1
X_11383_ _02246_ _03697_ _03699_ _02249_ VGND VGND VPWR VPWR _03726_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_34_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10755__A2 _01061_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10334_ _02372_ _02573_ VGND VGND VPWR VPWR _02574_ sky130_fd_sc_hd__nand2_1
X_13122_ _05637_ _05638_ VGND VGND VPWR VPWR _05639_ sky130_fd_sc_hd__nand2_1
XFILLER_0_131_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13053_ _05546_ _05562_ VGND VGND VPWR VPWR _05563_ sky130_fd_sc_hd__and2_2
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10265_ _00991_ _01356_ _01756_ _02294_ _02497_ VGND VGND VPWR VPWR _02498_ sky130_fd_sc_hd__a41oi_4
XANTENNA__10291__A _05577_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12004_ _00257_ _00670_ _02090_ _01780_ VGND VGND VPWR VPWR _04409_ sky130_fd_sc_hd__and4_1
X_10196_ _02082_ _02422_ VGND VGND VPWR VPWR _02424_ sky130_fd_sc_hd__xor2_2
XFILLER_0_108_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13955_ _06353_ _06536_ VGND VGND VPWR VPWR _06537_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12906_ _05248_ _05400_ VGND VGND VPWR VPWR _05402_ sky130_fd_sc_hd__nand2_1
XANTENNA__09304__B _01352_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13886_ _06442_ _06444_ VGND VGND VPWR VPWR _06462_ sky130_fd_sc_hd__and2_1
XFILLER_0_76_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07105__A _00508_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12837_ _02728_ _05100_ _05277_ _05278_ VGND VGND VPWR VPWR _05326_ sky130_fd_sc_hd__o2bb2ai_2
XTAP_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12768_ _05248_ _05249_ VGND VGND VPWR VPWR _05250_ sky130_fd_sc_hd__nand2_1
XANTENNA__11673__A1_N _06733_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07759__B _06885_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11719_ _00262_ _01585_ _04095_ VGND VGND VPWR VPWR _04096_ sky130_fd_sc_hd__and3_1
XFILLER_0_37_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12699_ _04926_ _05033_ VGND VGND VPWR VPWR _05174_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_127_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput10 a[18] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__buf_4
XFILLER_0_142_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput21 a[28] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_126_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput32 a[9] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__buf_2
Xinput43 b[19] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__buf_2
XFILLER_0_3_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput54 b[29] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_40_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08930_ _00690_ _00861_ _00865_ VGND VGND VPWR VPWR _01038_ sky130_fd_sc_hd__or3_1
XANTENNA__08723__A1_N _00508_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08861_ _01372_ net46 VGND VGND VPWR VPWR _00962_ sky130_fd_sc_hd__nand2_1
X_07812_ _00563_ _06818_ _06820_ _00639_ VGND VGND VPWR VPWR _06941_ sky130_fd_sc_hd__a22o_1
X_08792_ _00804_ _00885_ VGND VGND VPWR VPWR _00887_ sky130_fd_sc_hd__or2_1
XANTENNA__13448__A1 _01252_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13448__B2 _01182_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07743_ _06870_ _06871_ VGND VGND VPWR VPWR _06872_ sky130_fd_sc_hd__and2_1
XFILLER_0_74_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07674_ net36 VGND VGND VPWR VPWR _06744_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__07678__A2 _06765_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09413_ _01565_ VGND VGND VPWR VPWR _01566_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09344_ _01488_ _01489_ _01486_ VGND VGND VPWR VPWR _01490_ sky130_fd_sc_hd__or3b_1
XFILLER_0_48_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09275_ _01414_ VGND VGND VPWR VPWR _01415_ sky130_fd_sc_hd__buf_4
XFILLER_0_114_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_859 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08226_ _02116_ _00112_ _00268_ _02149_ VGND VGND VPWR VPWR _00270_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09588__C1 _01752_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08157_ _00194_ _00199_ _00200_ VGND VGND VPWR VPWR _00201_ sky130_fd_sc_hd__a21o_1
XFILLER_0_43_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13687__A _01288_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07108_ _00541_ _00300_ VGND VGND VPWR VPWR _00552_ sky130_fd_sc_hd__nand2_1
X_08088_ _00110_ _00130_ _00131_ _00128_ VGND VGND VPWR VPWR _00132_ sky130_fd_sc_hd__o22a_1
XFILLER_0_101_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10050_ _01855_ _02262_ VGND VGND VPWR VPWR _02264_ sky130_fd_sc_hd__or2_1
XANTENNA__11935__A _00003_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13740_ _05870_ _05873_ VGND VGND VPWR VPWR _06301_ sky130_fd_sc_hd__nor2_1
X_10952_ _03251_ _03252_ VGND VGND VPWR VPWR _03253_ sky130_fd_sc_hd__or2b_1
XFILLER_0_97_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13671_ _01183_ _02766_ _06223_ VGND VGND VPWR VPWR _06225_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_97_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10883_ _03135_ _03124_ _03134_ VGND VGND VPWR VPWR _03177_ sky130_fd_sc_hd__nor3_1
XFILLER_0_85_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08963__B _01076_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11670__A _07010_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12622_ _05041_ _05042_ _05084_ VGND VGND VPWR VPWR _05089_ sky130_fd_sc_hd__and3_1
XANTENNA__12485__B _00779_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12553_ _05004_ _05006_ _05009_ VGND VGND VPWR VPWR _05013_ sky130_fd_sc_hd__nand3_1
X_11504_ _03853_ _03857_ _03858_ VGND VGND VPWR VPWR _03859_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_41_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12484_ _00374_ _00741_ _04935_ _04936_ VGND VGND VPWR VPWR _04937_ sky130_fd_sc_hd__a31o_1
XFILLER_0_34_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14223_ _00406_ _00408_ VGND VGND VPWR VPWR _06807_ sky130_fd_sc_hd__and2_1
X_11435_ _03748_ VGND VGND VPWR VPWR _03783_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_110_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11366_ _03693_ _03695_ _03706_ VGND VGND VPWR VPWR _03708_ sky130_fd_sc_hd__o21a_1
X_14154_ _06619_ _06632_ _06635_ VGND VGND VPWR VPWR _06753_ sky130_fd_sc_hd__or3_2
X_13105_ _04028_ _05619_ VGND VGND VPWR VPWR _05620_ sky130_fd_sc_hd__xnor2_4
X_10317_ _02553_ _02555_ VGND VGND VPWR VPWR _02556_ sky130_fd_sc_hd__xnor2_1
X_14085_ _06102_ _06650_ _06676_ VGND VGND VPWR VPWR _06679_ sky130_fd_sc_hd__nor3_1
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11297_ _02810_ _02899_ _02901_ _03632_ VGND VGND VPWR VPWR _03633_ sky130_fd_sc_hd__a211o_1
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10452__C _02703_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10248_ _02391_ _02150_ _02479_ VGND VGND VPWR VPWR _02481_ sky130_fd_sc_hd__and3_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13036_ _05540_ _05542_ _05530_ VGND VGND VPWR VPWR _05545_ sky130_fd_sc_hd__a21o_1
XANTENNA__07357__A1 _01744_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10179_ _02403_ _03894_ _06744_ _02400_ VGND VGND VPWR VPWR _02405_ sky130_fd_sc_hd__and4b_1
XFILLER_0_28_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08857__C net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09315__A _00262_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13938_ _06514_ _06517_ VGND VGND VPWR VPWR _06519_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13869_ _06423_ _06430_ VGND VGND VPWR VPWR _06443_ sky130_fd_sc_hd__and2_1
XFILLER_0_147_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07390_ _02949_ _03631_ VGND VGND VPWR VPWR _03642_ sky130_fd_sc_hd__nand2_2
XANTENNA__13602__A1 _01061_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12395__B _00613_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09060_ _01179_ VGND VGND VPWR VPWR _01180_ sky130_fd_sc_hd__buf_4
XANTENNA__09985__A _06937_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08011_ _00053_ _00054_ VGND VGND VPWR VPWR _00055_ sky130_fd_sc_hd__or2_1
XFILLER_0_71_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09962_ _02165_ _02166_ VGND VGND VPWR VPWR _02167_ sky130_fd_sc_hd__xor2_2
XFILLER_0_100_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08913_ _00830_ _01017_ VGND VGND VPWR VPWR _01019_ sky130_fd_sc_hd__or2_1
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09893_ _06626_ _02090_ _02088_ _06450_ VGND VGND VPWR VPWR _02091_ sky130_fd_sc_hd__a22oi_1
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08844_ _00940_ _00942_ VGND VGND VPWR VPWR _00943_ sky130_fd_sc_hd__xnor2_4
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08775_ _00513_ _00520_ _00701_ VGND VGND VPWR VPWR _00868_ sky130_fd_sc_hd__o21a_1
XFILLER_0_79_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07726_ _06790_ _06850_ VGND VGND VPWR VPWR _06855_ sky130_fd_sc_hd__nand2_1
XANTENNA__10104__B1 _02158_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07657_ _06263_ _06549_ VGND VGND VPWR VPWR _06560_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12586__A _03707_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07588_ _03103_ _05800_ VGND VGND VPWR VPWR _05808_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09327_ _00145_ VGND VGND VPWR VPWR _01472_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_48_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10537__C _02724_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09258_ _01099_ _01395_ VGND VGND VPWR VPWR _01397_ sky130_fd_sc_hd__nor2_1
XFILLER_0_51_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08209_ _00081_ _00176_ _00100_ VGND VGND VPWR VPWR _00253_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_106_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09189_ _00257_ _00670_ _00819_ _00818_ VGND VGND VPWR VPWR _01321_ sky130_fd_sc_hd__nand4_1
XFILLER_0_50_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11220_ _03545_ _03546_ _03547_ VGND VGND VPWR VPWR _03548_ sky130_fd_sc_hd__a21o_1
XFILLER_0_43_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10553__B _02993_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11151_ _03244_ _03172_ VGND VGND VPWR VPWR _03472_ sky130_fd_sc_hd__nand2_1
X_10102_ _02318_ _02319_ VGND VGND VPWR VPWR _02320_ sky130_fd_sc_hd__or2_1
XFILLER_0_101_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11082_ _03394_ _03395_ VGND VGND VPWR VPWR _03396_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07339__A1 _03070_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07339__B2 _02280_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10033_ _01735_ _01851_ _01850_ VGND VGND VPWR VPWR _02245_ sky130_fd_sc_hd__o21ba_1
XANTENNA__11665__A _06885_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09135__A _05456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11984_ _04383_ _04384_ _04382_ VGND VGND VPWR VPWR _04387_ sky130_fd_sc_hd__a21o_1
XFILLER_0_86_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13723_ _06272_ _06278_ _06280_ VGND VGND VPWR VPWR _06282_ sky130_fd_sc_hd__or3_1
X_10935_ _02538_ _02540_ _03233_ VGND VGND VPWR VPWR _03234_ sky130_fd_sc_hd__a21o_1
XFILLER_0_85_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13654_ _06199_ _06205_ VGND VGND VPWR VPWR _06206_ sky130_fd_sc_hd__xnor2_1
X_10866_ _03156_ _03157_ VGND VGND VPWR VPWR _03159_ sky130_fd_sc_hd__and2_1
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12605_ _05068_ _05069_ VGND VGND VPWR VPWR _05070_ sky130_fd_sc_hd__nand2_1
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13585_ _06018_ _05985_ _06121_ _06129_ VGND VGND VPWR VPWR _06130_ sky130_fd_sc_hd__and4_1
XFILLER_0_137_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_859 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10797_ _03061_ _03060_ VGND VGND VPWR VPWR _03083_ sky130_fd_sc_hd__and2b_1
XPHY_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12536_ _04982_ _04984_ VGND VGND VPWR VPWR _04995_ sky130_fd_sc_hd__nand2_1
XFILLER_0_124_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13348__B1 _02305_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12467_ _04915_ _04918_ VGND VGND VPWR VPWR _04919_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_output92_A net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14206_ _02270_ _06796_ VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__xnor2_4
XFILLER_0_111_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11418_ _03739_ _03764_ VGND VGND VPWR VPWR _03765_ sky130_fd_sc_hd__or2_1
XANTENNA__11559__B _01960_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08214__A _00114_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12398_ _00374_ _01584_ VGND VGND VPWR VPWR _04843_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14137_ _06730_ _06734_ VGND VGND VPWR VPWR _06735_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11349_ _02249_ _01312_ _01956_ VGND VGND VPWR VPWR _03689_ sky130_fd_sc_hd__and3_1
XFILLER_0_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14068_ _06108_ _06079_ VGND VGND VPWR VPWR _06661_ sky130_fd_sc_hd__and2b_1
XANTENNA__11575__A _00263_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13019_ _01639_ _02046_ VGND VGND VPWR VPWR _05526_ sky130_fd_sc_hd__and2_1
X_08560_ _00542_ _00545_ VGND VGND VPWR VPWR _00633_ sky130_fd_sc_hd__and2b_1
X_07511_ _04345_ _04356_ _04829_ VGND VGND VPWR VPWR _04972_ sky130_fd_sc_hd__and3_1
XFILLER_0_76_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08491_ _00553_ _00557_ VGND VGND VPWR VPWR _00558_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_9_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07442_ _03587_ _04103_ _04191_ _03576_ VGND VGND VPWR VPWR _04213_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10638__B _02858_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07373_ _02839_ _03433_ _03444_ VGND VGND VPWR VPWR _03455_ sky130_fd_sc_hd__nor3_2
XFILLER_0_18_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13014__B _05494_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08108__B _00094_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09112_ _00943_ _01235_ _01236_ VGND VGND VPWR VPWR _01237_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_17_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10357__C _00423_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12853__B _01586_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09043_ _01115_ _01160_ VGND VGND VPWR VPWR _01161_ sky130_fd_sc_hd__xor2_1
XFILLER_0_5_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_328 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07947__B _07075_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09865__D _03740_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap140 _03455_ VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_102_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12562__A1 _00380_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09945_ _02145_ _02147_ VGND VGND VPWR VPWR _02148_ sky130_fd_sc_hd__xnor2_2
XANTENNA__09881__C _00413_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08778__B _00871_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09876_ _02070_ _02071_ VGND VGND VPWR VPWR _02073_ sky130_fd_sc_hd__xnor2_1
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08827_ _00901_ _03762_ _00753_ _00752_ VGND VGND VPWR VPWR _00925_ sky130_fd_sc_hd__a31o_1
XTAP_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08758_ _00848_ _00849_ VGND VGND VPWR VPWR _00850_ sky130_fd_sc_hd__nor2_1
XANTENNA__08794__A _00765_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07709_ _06832_ _06837_ VGND VGND VPWR VPWR _06838_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11932__B _01272_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08689_ _00602_ _00772_ VGND VGND VPWR VPWR _00774_ sky130_fd_sc_hd__nor2_1
XANTENNA__10829__A _01350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10720_ _02990_ _02995_ _02997_ VGND VGND VPWR VPWR _02998_ sky130_fd_sc_hd__a21oi_1
XTAP_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09246__A1 _03268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10651_ _02891_ _02881_ VGND VGND VPWR VPWR _02922_ sky130_fd_sc_hd__or2b_1
XFILLER_0_82_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09246__B2 _05577_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07257__B1 _00333_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10582_ _00310_ _01413_ VGND VGND VPWR VPWR _02846_ sky130_fd_sc_hd__nand2_1
X_13370_ _05891_ _05894_ VGND VGND VPWR VPWR _05895_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09797__A2 _01585_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12321_ _04744_ _04757_ VGND VGND VPWR VPWR _04758_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_188 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12252_ _00378_ _02120_ VGND VGND VPWR VPWR _04682_ sky130_fd_sc_hd__nand2_1
XANTENNA__08757__B1 _00846_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11203_ _03500_ _03502_ _03503_ _03501_ VGND VGND VPWR VPWR _03529_ sky130_fd_sc_hd__o22a_1
X_12183_ _02382_ _02385_ _02588_ _04603_ _04605_ VGND VGND VPWR VPWR _04606_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_102_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11134_ _03450_ _03452_ VGND VGND VPWR VPWR _03453_ sky130_fd_sc_hd__and2_2
XFILLER_0_102_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07592__B _05588_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11065_ _03363_ _03376_ VGND VGND VPWR VPWR _03377_ sky130_fd_sc_hd__nor2_1
X_10016_ _02223_ _02225_ VGND VGND VPWR VPWR _02227_ sky130_fd_sc_hd__nand2_1
XANTENNA__09182__B1 _00526_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11967_ _04296_ net144 _04368_ VGND VGND VPWR VPWR _04369_ sky130_fd_sc_hd__o21a_1
XFILLER_0_58_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08288__A2 _00094_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13706_ _01288_ _02720_ _02725_ _00416_ VGND VGND VPWR VPWR _06264_ sky130_fd_sc_hd__a22o_1
X_10918_ _03212_ _03214_ VGND VGND VPWR VPWR _03216_ sky130_fd_sc_hd__and2_1
X_11898_ _06428_ _01954_ _02135_ _06439_ VGND VGND VPWR VPWR _04293_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_117_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13637_ _06185_ _06187_ VGND VGND VPWR VPWR _06188_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10849_ _05742_ _00541_ _01545_ net52 VGND VGND VPWR VPWR _03140_ sky130_fd_sc_hd__and4_1
XANTENNA__10177__C _03685_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13568_ _06102_ _06103_ _06110_ VGND VGND VPWR VPWR _06112_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09966__C net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12792__A1 _00392_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12792__B2 _00389_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12519_ _04958_ _04965_ _04966_ VGND VGND VPWR VPWR _04976_ sky130_fd_sc_hd__o21a_1
XANTENNA__10474__A net57 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13499_ _06009_ _06018_ _03687_ _03684_ VGND VGND VPWR VPWR _06036_ sky130_fd_sc_hd__and4_1
XFILLER_0_2_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_394 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07783__A _01044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07991_ _07030_ _00034_ VGND VGND VPWR VPWR _00035_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09730_ _01686_ _01688_ VGND VGND VPWR VPWR _01913_ sky130_fd_sc_hd__or2b_1
X_09661_ _01649_ _01837_ VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__xor2_4
X_08612_ _06428_ _06439_ _00144_ _00298_ VGND VGND VPWR VPWR _00690_ sky130_fd_sc_hd__and4_1
X_09592_ _06818_ net8 net9 _06820_ VGND VGND VPWR VPWR _01762_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09503__A _01508_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08543_ _01230_ _00612_ _00613_ _01284_ VGND VGND VPWR VPWR _00614_ sky130_fd_sc_hd__a22o_1
XANTENNA__11871__A2_N _01601_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08474_ _00528_ _00529_ _00537_ VGND VGND VPWR VPWR _00539_ sky130_fd_sc_hd__nor3_1
XFILLER_0_119_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_455 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07425_ _04015_ VGND VGND VPWR VPWR _04026_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_119_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07356_ _02719_ VGND VGND VPWR VPWR _03268_ sky130_fd_sc_hd__buf_4
XFILLER_0_73_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12583__B _01412_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_188 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07287_ _01098_ _01142_ VGND VGND VPWR VPWR _02510_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09026_ _01134_ _01141_ VGND VGND VPWR VPWR _01143_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_372 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13695__A _02426_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07693__A _00891_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07411__B1 _03718_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09951__A2 _01410_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09928_ _02112_ _02113_ _02129_ VGND VGND VPWR VPWR _02130_ sky130_fd_sc_hd__a21o_1
XANTENNA__12838__A2 _02724_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09859_ _01868_ _01950_ VGND VGND VPWR VPWR _02054_ sky130_fd_sc_hd__nor2_1
X_12870_ _05360_ _05361_ VGND VGND VPWR VPWR _05362_ sky130_fd_sc_hd__nand2_1
XTAP_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11662__B _06765_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11821_ _04203_ _04204_ _04207_ VGND VGND VPWR VPWR _04208_ sky130_fd_sc_hd__o21a_1
XTAP_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11752_ _02615_ _04128_ _04130_ VGND VGND VPWR VPWR _04132_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_56_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_455 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10703_ _00388_ _03004_ _01059_ _01412_ VGND VGND VPWR VPWR _02979_ sky130_fd_sc_hd__and4_1
XTAP_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14212__A1 _00464_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11683_ _04041_ _04046_ VGND VGND VPWR VPWR _04056_ sky130_fd_sc_hd__xnor2_1
XTAP_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14212__B2 _02051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13422_ _05949_ _05951_ VGND VGND VPWR VPWR _05952_ sky130_fd_sc_hd__and2_1
X_10634_ _02901_ _02902_ VGND VGND VPWR VPWR _02903_ sky130_fd_sc_hd__nor2_1
XANTENNA__12223__B1 _02117_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13353_ _05341_ _05347_ VGND VGND VPWR VPWR _05876_ sky130_fd_sc_hd__and2_1
XFILLER_0_23_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10294__A _03268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10565_ _02804_ _02801_ VGND VGND VPWR VPWR _02827_ sky130_fd_sc_hd__or2b_1
XFILLER_0_63_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12304_ _04737_ _04738_ _00608_ _01601_ VGND VGND VPWR VPWR _04739_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_106_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13284_ _05725_ _05806_ VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__xnor2_1
X_10496_ _00636_ _00526_ _02735_ _02731_ VGND VGND VPWR VPWR _02752_ sky130_fd_sc_hd__and4_1
XFILLER_0_122_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12235_ _00783_ _00778_ _01178_ _01248_ VGND VGND VPWR VPWR _04663_ sky130_fd_sc_hd__and4_1
XANTENNA__08699__A _01383_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12166_ _04519_ _04530_ VGND VGND VPWR VPWR _04588_ sky130_fd_sc_hd__and2_1
X_11117_ _03428_ _03427_ VGND VGND VPWR VPWR _03435_ sky130_fd_sc_hd__or2_1
X_12097_ _04374_ _04380_ _04441_ VGND VGND VPWR VPWR _04512_ sky130_fd_sc_hd__o21a_1
XANTENNA__07108__A _00541_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11048_ _03346_ _03349_ _03350_ VGND VGND VPWR VPWR _03359_ sky130_fd_sc_hd__a21oi_1
Xinput8 a[16] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_127_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10469__A _02721_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12999_ _05487_ _05503_ VGND VGND VPWR VPWR _05504_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_87_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07210_ _01613_ _01580_ VGND VGND VPWR VPWR _01667_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_129_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08190_ _00210_ _00214_ VGND VGND VPWR VPWR _00234_ sky130_fd_sc_hd__nand2_1
XANTENNA__12214__B1 _01254_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11902__A1_N _03070_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07141_ _00891_ _00901_ VGND VGND VPWR VPWR _00912_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10776__B1 _02727_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08402__A _00459_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07974_ _06961_ _07017_ _00017_ VGND VGND VPWR VPWR _00018_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09146__B1 _01211_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09713_ _01893_ VGND VGND VPWR VPWR _01894_ sky130_fd_sc_hd__inv_2
X_09644_ _01255_ _01571_ _01817_ VGND VGND VPWR VPWR _01819_ sky130_fd_sc_hd__o21a_1
XANTENNA__09233__A _00959_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09575_ _01738_ _01742_ VGND VGND VPWR VPWR _01743_ sky130_fd_sc_hd__nand2_1
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11913__D _03679_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08526_ _00570_ _00594_ VGND VGND VPWR VPWR _00596_ sky130_fd_sc_hd__or2_4
XANTENNA__10098__B net53 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08457_ _00516_ _00518_ VGND VGND VPWR VPWR _00521_ sky130_fd_sc_hd__and2_1
XFILLER_0_108_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07408_ _03751_ _03828_ VGND VGND VPWR VPWR _03839_ sky130_fd_sc_hd__nand2_1
X_08388_ _00978_ _00880_ _04180_ net43 VGND VGND VPWR VPWR _00445_ sky130_fd_sc_hd__and4_1
XFILLER_0_18_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07339_ _03070_ _02259_ _02171_ _02280_ VGND VGND VPWR VPWR _03081_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07838__D _06966_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11003__A _05192_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_823 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10350_ _02496_ _02498_ _02591_ VGND VGND VPWR VPWR _02592_ sky130_fd_sc_hd__a21o_1
XFILLER_0_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09009_ _03004_ _00113_ _00114_ _00094_ VGND VGND VPWR VPWR _01124_ sky130_fd_sc_hd__and4_1
XFILLER_0_130_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10281_ _02512_ _02515_ VGND VGND VPWR VPWR _02516_ sky130_fd_sc_hd__xor2_1
XFILLER_0_103_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12020_ _04425_ _04426_ VGND VGND VPWR VPWR _04427_ sky130_fd_sc_hd__xnor2_2
XANTENNA__08669__D net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13971_ _06541_ _06554_ VGND VGND VPWR VPWR _06555_ sky130_fd_sc_hd__and2_1
XANTENNA__08966__B net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12922_ _05417_ _05418_ VGND VGND VPWR VPWR _05419_ sky130_fd_sc_hd__nor2_1
XANTENNA__12488__B _00914_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11392__B _00268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12853_ _00572_ _01586_ _02306_ _02305_ VGND VGND VPWR VPWR _05343_ sky130_fd_sc_hd__and4_1
XTAP_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11804_ _04186_ _02677_ _04187_ VGND VGND VPWR VPWR _04189_ sky130_fd_sc_hd__a21o_1
XTAP_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12784_ _00414_ _00572_ _01411_ _02849_ VGND VGND VPWR VPWR _05267_ sky130_fd_sc_hd__and4_1
XTAP_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12995__A1 _00381_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11735_ _04109_ _04112_ VGND VGND VPWR VPWR _04113_ sky130_fd_sc_hd__nor2_1
XFILLER_0_113_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11666_ _04035_ _04036_ VGND VGND VPWR VPWR _04038_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_83_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13405_ _01066_ _03414_ _01955_ _03686_ VGND VGND VPWR VPWR _05933_ sky130_fd_sc_hd__and4_1
X_10617_ _02868_ _02884_ VGND VGND VPWR VPWR _02885_ sky130_fd_sc_hd__nor2_1
XFILLER_0_107_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11597_ _03940_ _03912_ _03936_ VGND VGND VPWR VPWR _03962_ sky130_fd_sc_hd__and3_1
XFILLER_0_3_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13336_ _00914_ _00745_ _02724_ _02728_ VGND VGND VPWR VPWR _05858_ sky130_fd_sc_hd__nand4_1
X_10548_ _00818_ _02725_ _02730_ _00819_ VGND VGND VPWR VPWR _02809_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13267_ _02495_ _05763_ _05788_ _05791_ VGND VGND VPWR VPWR _05792_ sky130_fd_sc_hd__a31o_4
XFILLER_0_122_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10479_ _01472_ _00636_ _02726_ _02730_ VGND VGND VPWR VPWR _02733_ sky130_fd_sc_hd__and4_1
XFILLER_0_110_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12218_ _04641_ _04644_ VGND VGND VPWR VPWR _04645_ sky130_fd_sc_hd__or2_1
XANTENNA__09915__A2 _01960_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11567__B _00497_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13198_ _05717_ _05718_ VGND VGND VPWR VPWR _05723_ sky130_fd_sc_hd__nor2_1
X_12149_ _04558_ _04561_ _04559_ VGND VGND VPWR VPWR _04569_ sky130_fd_sc_hd__or3_1
XFILLER_0_47_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12679__A _05136_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07690_ _06818_ VGND VGND VPWR VPWR _06819_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08351__A1 _00464_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07154__A2 _01044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12398__B _01584_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10199__A _02090_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09360_ _01507_ VGND VGND VPWR VPWR _01508_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_93_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08892__A _03543_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08311_ _06998_ _06999_ VGND VGND VPWR VPWR _00361_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_74_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09291_ _01243_ _01432_ VGND VGND VPWR VPWR _01433_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_47_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08242_ _00283_ _00284_ VGND VGND VPWR VPWR _00286_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07301__A net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_423 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08173_ _06120_ _00212_ VGND VGND VPWR VPWR _00217_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_144_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09603__A1 _06428_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08116__B _00142_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09603__B2 _06439_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07124_ net27 _00705_ net28 net161 VGND VGND VPWR VPWR _00726_ sky130_fd_sc_hd__and4_1
XFILLER_0_125_491 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07955__B _00497_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput120 net120 VGND VGND VPWR VPWR prod[5] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_30_459 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12580__C _02849_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09228__A _04048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07917__A1 net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07917__B2 net61 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07957_ _03554_ _00410_ _03015_ _00519_ VGND VGND VPWR VPWR _00001_ sky130_fd_sc_hd__a22o_1
X_07888_ _07008_ _07016_ VGND VGND VPWR VPWR _07017_ sky130_fd_sc_hd__xor2_1
XANTENNA__08906__A1_N _00003_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09627_ _01796_ _01800_ VGND VGND VPWR VPWR _01801_ sky130_fd_sc_hd__and2b_1
XFILLER_0_97_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09558_ _00844_ _00635_ _07040_ _00843_ VGND VGND VPWR VPWR _01725_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_38_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08509_ _01744_ _00311_ _00413_ _00571_ VGND VGND VPWR VPWR _00577_ sky130_fd_sc_hd__and4_1
XFILLER_0_136_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09489_ _01647_ _01648_ VGND VGND VPWR VPWR _01649_ sky130_fd_sc_hd__nand2_2
XFILLER_0_65_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11520_ _03869_ _03876_ VGND VGND VPWR VPWR _03877_ sky130_fd_sc_hd__xor2_4
XFILLER_0_135_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11451_ _06964_ _00121_ _01953_ _02133_ VGND VGND VPWR VPWR _03801_ sky130_fd_sc_hd__and4_1
XFILLER_0_61_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10402_ _05445_ _01177_ _01247_ _05467_ VGND VGND VPWR VPWR _02649_ sky130_fd_sc_hd__a22o_1
X_14170_ _06768_ _06769_ VGND VGND VPWR VPWR _06770_ sky130_fd_sc_hd__and2b_1
X_11382_ _02246_ _02249_ _03697_ _03699_ VGND VGND VPWR VPWR _03725_ sky130_fd_sc_hd__and4_1
XFILLER_0_104_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13121_ _05608_ _05620_ VGND VGND VPWR VPWR _05638_ sky130_fd_sc_hd__xor2_2
XFILLER_0_0_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10333_ _02569_ _02572_ VGND VGND VPWR VPWR _02573_ sky130_fd_sc_hd__xor2_1
XFILLER_0_131_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13052_ _05548_ _05561_ VGND VGND VPWR VPWR _05562_ sky130_fd_sc_hd__xnor2_4
X_10264_ _01757_ _02294_ VGND VGND VPWR VPWR _02497_ sky130_fd_sc_hd__and2_1
XANTENNA__07584__C _00901_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08042__A _00002_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10291__B _01410_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12003_ _04340_ _04342_ VGND VGND VPWR VPWR _04408_ sky130_fd_sc_hd__and2b_1
X_10195_ _02392_ _02421_ VGND VGND VPWR VPWR _02422_ sky130_fd_sc_hd__xor2_2
XANTENNA__07881__A net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13954_ _06354_ _06343_ VGND VGND VPWR VPWR _06536_ sky130_fd_sc_hd__and2b_1
XFILLER_0_17_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12905_ _05232_ _05249_ VGND VGND VPWR VPWR _05400_ sky130_fd_sc_hd__nand2_1
X_13885_ _06454_ _06455_ _06459_ VGND VGND VPWR VPWR _06460_ sky130_fd_sc_hd__o21ai_2
XANTENNA__10140__A1 _00458_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_459 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12836_ _05279_ _05322_ _05323_ VGND VGND VPWR VPWR _05325_ sky130_fd_sc_hd__a21o_1
XTAP_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12767_ _04654_ _04659_ _05246_ _05245_ VGND VGND VPWR VPWR _05249_ sky130_fd_sc_hd__a31o_1
XFILLER_0_29_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14219__A _06804_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09833__A1 _07004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09320__B _01463_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11718_ _00263_ _01600_ VGND VGND VPWR VPWR _04095_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_222 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12698_ _05167_ _05172_ VGND VGND VPWR VPWR _05173_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_140_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput11 a[19] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_4
X_11649_ _03708_ _03731_ _03733_ VGND VGND VPWR VPWR _04019_ sky130_fd_sc_hd__a21o_1
Xinput22 a[29] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_71_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput33 b[0] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__buf_6
Xinput44 b[1] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_3_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput55 b[2] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__buf_6
XFILLER_0_107_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13319_ _05792_ _05807_ _05836_ _05838_ _05840_ VGND VGND VPWR VPWR _05841_ sky130_fd_sc_hd__a311o_4
XANTENNA__10482__A _02735_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08860_ _00958_ _00960_ VGND VGND VPWR VPWR _00961_ sky130_fd_sc_hd__or2b_1
X_07811_ net27 net28 _06818_ net34 VGND VGND VPWR VPWR _06940_ sky130_fd_sc_hd__and4_1
X_08791_ _00804_ _00885_ VGND VGND VPWR VPWR _00886_ sky130_fd_sc_hd__and2_1
XANTENNA__13448__A2 _02736_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07742_ _06755_ _06869_ VGND VGND VPWR VPWR _06871_ sky130_fd_sc_hd__or2_1
X_07673_ net37 VGND VGND VPWR VPWR _06733_ sky130_fd_sc_hd__clkbuf_4
X_09412_ _04510_ _01177_ _01246_ _00661_ VGND VGND VPWR VPWR _01565_ sky130_fd_sc_hd__a22o_1
XANTENNA__08262__A1_N _03059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09343_ _00557_ _01167_ _01441_ _01442_ VGND VGND VPWR VPWR _01489_ sky130_fd_sc_hd__a31o_1
XANTENNA__13081__B1 _05593_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11631__A1 _01155_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09274_ _01413_ VGND VGND VPWR VPWR _01414_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_90_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08225_ _02116_ _02149_ _00112_ _00268_ VGND VGND VPWR VPWR _00269_ sky130_fd_sc_hd__and4_1
XFILLER_0_74_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_214 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08156_ _00196_ _00198_ VGND VGND VPWR VPWR _00200_ sky130_fd_sc_hd__nor2_1
XANTENNA__13687__B _02090_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07107_ net29 VGND VGND VPWR VPWR _00541_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_30_223 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08260__B1 _04928_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08087_ _00032_ _00127_ _00110_ VGND VGND VPWR VPWR _00131_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_101_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11935__B _01585_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08989_ _01068_ _01069_ _01101_ VGND VGND VPWR VPWR _01102_ sky130_fd_sc_hd__o21a_1
XFILLER_0_98_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10951_ _00143_ _01508_ _01505_ _04906_ VGND VGND VPWR VPWR _03252_ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_407 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13670_ _01183_ _06074_ _06223_ VGND VGND VPWR VPWR _06224_ sky130_fd_sc_hd__nand3_1
X_10882_ _03093_ _03175_ VGND VGND VPWR VPWR _03176_ sky130_fd_sc_hd__nor2_1
XANTENNA__08963__C net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11670__B net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09421__A _00138_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12621_ _05086_ _05087_ VGND VGND VPWR VPWR _05088_ sky130_fd_sc_hd__or2_2
XANTENNA__12485__C _00742_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11622__A1 _00519_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12552_ _04865_ _05011_ VGND VGND VPWR VPWR _05012_ sky130_fd_sc_hd__nor2_2
XFILLER_0_136_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11503_ _03840_ _03842_ VGND VGND VPWR VPWR _03858_ sky130_fd_sc_hd__xor2_1
XFILLER_0_81_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12483_ _00612_ _00777_ _00423_ _03762_ VGND VGND VPWR VPWR _04936_ sky130_fd_sc_hd__and4_1
XANTENNA__12782__A _01600_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_359 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14222_ _00401_ _06806_ VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__xnor2_2
X_11434_ _03780_ _03781_ VGND VGND VPWR VPWR _03782_ sky130_fd_sc_hd__or2b_1
XANTENNA__07876__A _02467_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14153_ _06750_ _06751_ VGND VGND VPWR VPWR _06752_ sky130_fd_sc_hd__nand2_2
X_11365_ _03704_ _03705_ VGND VGND VPWR VPWR _03706_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_22_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13104_ _05609_ _05615_ _05617_ _05618_ VGND VGND VPWR VPWR _05619_ sky130_fd_sc_hd__o31a_2
XFILLER_0_0_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10316_ _04598_ net45 VGND VGND VPWR VPWR _02555_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14084_ _06677_ VGND VGND VPWR VPWR _06678_ sky130_fd_sc_hd__inv_2
X_11296_ _00819_ _00818_ _02736_ _02737_ VGND VGND VPWR VPWR _03632_ sky130_fd_sc_hd__and4_1
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13035_ _05530_ _05540_ _05542_ VGND VGND VPWR VPWR _05543_ sky130_fd_sc_hd__and3_1
X_10247_ _02391_ _02150_ _02479_ VGND VGND VPWR VPWR _02480_ sky130_fd_sc_hd__a21oi_2
XANTENNA__07357__A2 _03268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10178_ _06744_ _03773_ _02402_ _02403_ VGND VGND VPWR VPWR _02404_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__08857__D net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09315__B _00859_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12022__A _06626_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07116__A net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13937_ _06514_ _06517_ VGND VGND VPWR VPWR _06518_ sky130_fd_sc_hd__nor2_1
XFILLER_0_135_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13868_ _06438_ _06441_ VGND VGND VPWR VPWR _06442_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12819_ _05304_ _05305_ VGND VGND VPWR VPWR _05306_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10477__A _02730_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13799_ _02187_ _02189_ _03686_ _03683_ VGND VGND VPWR VPWR _06366_ sky130_fd_sc_hd__and4_1
XFILLER_0_56_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13602__A2 _03783_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12395__C _00413_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09985__B _06637_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08010_ _00047_ _00052_ VGND VGND VPWR VPWR _00054_ sky130_fd_sc_hd__and2_1
XANTENNA__07786__A _01000_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09961_ _01661_ _01929_ _01928_ VGND VGND VPWR VPWR _02166_ sky130_fd_sc_hd__a21o_1
XFILLER_0_40_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09560__A1_N _00654_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08912_ _00830_ _01017_ VGND VGND VPWR VPWR _01018_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09892_ _01601_ VGND VGND VPWR VPWR _02090_ sky130_fd_sc_hd__clkbuf_4
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08843_ _00596_ _00764_ _00941_ VGND VGND VPWR VPWR _00942_ sky130_fd_sc_hd__o21ai_4
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08774_ _00702_ VGND VGND VPWR VPWR _00867_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13970__B _06540_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07725_ _06852_ _06853_ VGND VGND VPWR VPWR _06854_ sky130_fd_sc_hd__or2_1
XANTENNA__10104__A1 _00650_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10104__B2 _02105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07656_ _06527_ _06538_ VGND VGND VPWR VPWR _06549_ sky130_fd_sc_hd__nor2_1
XANTENNA__12586__B _03740_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07587_ _05771_ _05790_ VGND VGND VPWR VPWR _05800_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09326_ _00526_ _01468_ _01469_ VGND VGND VPWR VPWR _01471_ sky130_fd_sc_hd__a21bo_1
XANTENNA__10188__A2_N _00734_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09257_ _01099_ _01395_ VGND VGND VPWR VPWR _01396_ sky130_fd_sc_hd__and2_1
XANTENNA__10537__D _02728_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08208_ _00081_ _00176_ VGND VGND VPWR VPWR _00252_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09188_ _00257_ _00293_ _00294_ _00670_ VGND VGND VPWR VPWR _01320_ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08139_ _00089_ _00090_ _00182_ VGND VGND VPWR VPWR _00183_ sky130_fd_sc_hd__and3_1
XFILLER_0_120_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10553__C _02168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11011__A _04598_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11150_ _03459_ _03460_ VGND VGND VPWR VPWR _03471_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_101_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10101_ _01934_ _02172_ _02317_ VGND VGND VPWR VPWR _02319_ sky130_fd_sc_hd__a21oi_1
X_11081_ _03375_ _03377_ VGND VGND VPWR VPWR _03395_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07339__A2 _02259_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10032_ _01489_ _01488_ _02243_ _01867_ VGND VGND VPWR VPWR _02244_ sky130_fd_sc_hd__o211a_2
XANTENNA__11665__B _01601_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09135__B _05478_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11983_ _04354_ _04355_ _04353_ VGND VGND VPWR VPWR _04386_ sky130_fd_sc_hd__a21o_1
X_13722_ _06272_ _06278_ _06280_ VGND VGND VPWR VPWR _06281_ sky130_fd_sc_hd__o21ai_1
X_10934_ _02504_ _02537_ VGND VGND VPWR VPWR _03233_ sky130_fd_sc_hd__and2b_1
XFILLER_0_86_727 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13653_ _06204_ _06196_ VGND VGND VPWR VPWR _06205_ sky130_fd_sc_hd__nor2_1
X_10865_ _03149_ _03152_ VGND VGND VPWR VPWR _03157_ sky130_fd_sc_hd__xor2_1
X_12604_ _05064_ _05061_ VGND VGND VPWR VPWR _05069_ sky130_fd_sc_hd__xnor2_1
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13584_ _06126_ _06127_ _06128_ VGND VGND VPWR VPWR _06129_ sky130_fd_sc_hd__and3_1
XFILLER_0_38_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10796_ _03079_ _03080_ VGND VGND VPWR VPWR _03082_ sky130_fd_sc_hd__nand2_1
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12535_ _04930_ _04992_ VGND VGND VPWR VPWR _04993_ sky130_fd_sc_hd__xor2_2
XFILLER_0_121_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13348__A1 _01584_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13348__B2 _01586_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12466_ _04869_ _04916_ VGND VGND VPWR VPWR _04918_ sky130_fd_sc_hd__nor2_1
XFILLER_0_124_567 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14205_ _02346_ _06795_ VGND VGND VPWR VPWR _06796_ sky130_fd_sc_hd__nand2_2
XFILLER_0_50_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13120__B _05636_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11417_ _00003_ _03738_ _03736_ _03737_ VGND VGND VPWR VPWR _03764_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_105_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12397_ _04830_ _04828_ VGND VGND VPWR VPWR _04842_ sky130_fd_sc_hd__and2b_1
X_14136_ _06731_ _06732_ VGND VGND VPWR VPWR _06734_ sky130_fd_sc_hd__nand2_1
X_11348_ _02249_ _01956_ _03687_ _01312_ VGND VGND VPWR VPWR _03688_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_773 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14067_ _06657_ _06659_ VGND VGND VPWR VPWR _06660_ sky130_fd_sc_hd__nand2_1
X_11279_ _03498_ _03511_ VGND VGND VPWR VPWR _03613_ sky130_fd_sc_hd__xor2_4
XANTENNA__09971__D _01411_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13018_ _05492_ _05507_ _05524_ VGND VGND VPWR VPWR _05525_ sky130_fd_sc_hd__and3_1
XANTENNA__11575__B _03750_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_705 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07510_ _04884_ _04950_ VGND VGND VPWR VPWR _04961_ sky130_fd_sc_hd__nand2_2
X_08490_ _00367_ _00554_ _00556_ VGND VGND VPWR VPWR _00557_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_89_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09061__A _01180_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07441_ _00431_ _04169_ _04180_ _04191_ VGND VGND VPWR VPWR _04202_ sky130_fd_sc_hd__and4_1
XFILLER_0_119_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07372_ _02456_ _02467_ _02861_ VGND VGND VPWR VPWR _03444_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_29_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_186 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09111_ _00984_ _01048_ VGND VGND VPWR VPWR _01236_ sky130_fd_sc_hd__and2_1
XFILLER_0_57_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09042_ _01116_ _01159_ VGND VGND VPWR VPWR _01160_ sky130_fd_sc_hd__xnor2_2
XANTENNA__12853__C _02306_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_142_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap130 _05595_ VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__clkbuf_2
Xmax_cap141 _06150_ VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__clkbuf_1
XANTENNA__12562__A2 _02008_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09944_ _02006_ _02028_ _02146_ VGND VGND VPWR VPWR _02147_ sky130_fd_sc_hd__o21a_1
XANTENNA__10670__A _00094_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09881__D _00572_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09875_ _01771_ _02022_ _02021_ VGND VGND VPWR VPWR _02071_ sky130_fd_sc_hd__a21o_1
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08826_ _00921_ _00922_ VGND VGND VPWR VPWR _00924_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08757_ _00669_ _00674_ _00846_ VGND VGND VPWR VPWR _00849_ sky130_fd_sc_hd__a21oi_1
XTAP_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07708_ net26 net63 VGND VGND VPWR VPWR _06837_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08688_ _00602_ _00772_ VGND VGND VPWR VPWR _00773_ sky130_fd_sc_hd__and2_1
XTAP_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10829__B _02728_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07639_ _06340_ _06351_ VGND VGND VPWR VPWR _06362_ sky130_fd_sc_hd__or2_1
XTAP_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13578__A1 _01250_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10650_ _02830_ _02838_ VGND VGND VPWR VPWR _02921_ sky130_fd_sc_hd__xor2_1
XANTENNA__09246__A2 _00612_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07257__A1 _02116_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09309_ _00843_ _00818_ _01451_ VGND VGND VPWR VPWR _01452_ sky130_fd_sc_hd__and3_1
XFILLER_0_75_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__07257__B2 _02171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10581_ _02843_ _02844_ VGND VGND VPWR VPWR _02845_ sky130_fd_sc_hd__or2b_1
XFILLER_0_146_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_679 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12320_ _04737_ _04739_ _04743_ VGND VGND VPWR VPWR _04757_ sky130_fd_sc_hd__nor3_1
XFILLER_0_90_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12251_ _04679_ _04680_ VGND VGND VPWR VPWR _04681_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_32_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08034__B _07075_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10013__B1 _00608_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11202_ _03523_ _03527_ VGND VGND VPWR VPWR _03528_ sky130_fd_sc_hd__nand2_1
XFILLER_0_121_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12182_ _03550_ _04604_ VGND VGND VPWR VPWR _04605_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10564__A1 _00818_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11133_ _03050_ _03451_ VGND VGND VPWR VPWR _03452_ sky130_fd_sc_hd__and2_1
XANTENNA__11676__A _00112_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11064_ _03362_ _03351_ _03361_ VGND VGND VPWR VPWR _03376_ sky130_fd_sc_hd__nor3_1
XANTENNA__08050__A _05203_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09182__A1 _00544_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10015_ _00459_ _02224_ VGND VGND VPWR VPWR _02225_ sky130_fd_sc_hd__nand2_1
XANTENNA__09182__B2 _01312_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13266__B1 _05789_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11966_ _04365_ _04366_ VGND VGND VPWR VPWR _04368_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12300__A _02190_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_604 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10917_ _03212_ _03214_ VGND VGND VPWR VPWR _03215_ sky130_fd_sc_hd__nor2_1
X_13705_ _06259_ _06261_ VGND VGND VPWR VPWR _06262_ sky130_fd_sc_hd__and2b_1
XFILLER_0_58_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11897_ _06417_ _06439_ _01954_ _02135_ VGND VGND VPWR VPWR _04292_ sky130_fd_sc_hd__and4_1
XFILLER_0_132_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13636_ _06184_ _06180_ VGND VGND VPWR VPWR _06187_ sky130_fd_sc_hd__and2b_1
XFILLER_0_39_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10848_ _00541_ _01545_ net52 _05742_ VGND VGND VPWR VPWR _03139_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10177__D _00423_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13567_ _06103_ _06110_ VGND VGND VPWR VPWR _06111_ sky130_fd_sc_hd__or2_1
XFILLER_0_125_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10779_ _03058_ _03062_ VGND VGND VPWR VPWR _03063_ sky130_fd_sc_hd__or2b_1
XFILLER_0_54_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08996__A1 _00464_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12518_ _04973_ _04974_ VGND VGND VPWR VPWR _04975_ sky130_fd_sc_hd__and2_1
XANTENNA__12792__A2 _02723_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13498_ _06018_ _03690_ _06034_ VGND VGND VPWR VPWR _06035_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_42_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08225__A _02116_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12449_ _04823_ _04811_ _04821_ VGND VGND VPWR VPWR _04899_ sky130_fd_sc_hd__and3_1
XFILLER_0_22_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10004__B1 _00613_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14119_ _06714_ _06715_ VGND VGND VPWR VPWR _06716_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07990_ _00032_ _00033_ VGND VGND VPWR VPWR _00034_ sky130_fd_sc_hd__and2_1
XANTENNA__10490__A _02247_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09660_ _01835_ _01836_ VGND VGND VPWR VPWR _01837_ sky130_fd_sc_hd__and2_2
X_08611_ _06428_ _00144_ _00310_ _06450_ VGND VGND VPWR VPWR _00689_ sky130_fd_sc_hd__a22oi_1
X_09591_ _06818_ _06820_ net9 VGND VGND VPWR VPWR _01761_ sky130_fd_sc_hd__and3_1
X_08542_ _04191_ VGND VGND VPWR VPWR _00613_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08473_ _00528_ _00529_ _00537_ VGND VGND VPWR VPWR _00538_ sky130_fd_sc_hd__o21a_1
XFILLER_0_147_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07424_ net41 VGND VGND VPWR VPWR _04015_ sky130_fd_sc_hd__buf_2
XFILLER_0_147_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07355_ _02675_ net189 VGND VGND VPWR VPWR _03257_ sky130_fd_sc_hd__nand2_1
XFILLER_0_116_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07286_ _01131_ _01109_ VGND VGND VPWR VPWR _02499_ sky130_fd_sc_hd__or2b_1
XFILLER_0_72_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09025_ _01139_ _01140_ VGND VGND VPWR VPWR _01141_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12880__A _00605_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13695__B _02737_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10546__A1 _00818_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07693__B _01120_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07411__B2 _01306_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09927_ _02126_ _02128_ VGND VGND VPWR VPWR _02129_ sky130_fd_sc_hd__xnor2_1
X_09858_ _01868_ _01950_ VGND VGND VPWR VPWR _02053_ sky130_fd_sc_hd__nand2_1
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08809_ _00903_ _00904_ VGND VGND VPWR VPWR _00905_ sky130_fd_sc_hd__xnor2_1
X_09789_ _02456_ _01181_ _01976_ VGND VGND VPWR VPWR _01978_ sky130_fd_sc_hd__a21o_1
XTAP_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11820_ _04182_ _04206_ VGND VGND VPWR VPWR _04207_ sky130_fd_sc_hd__xor2_1
XTAP_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11662__C _00414_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11751_ _02615_ _04128_ _04130_ VGND VGND VPWR VPWR _04131_ sky130_fd_sc_hd__and3_1
XTAP_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07478__B2 net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10702_ _02976_ _02977_ VGND VGND VPWR VPWR _02978_ sky130_fd_sc_hd__xnor2_1
XTAP_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11682_ _02606_ _02605_ VGND VGND VPWR VPWR _04055_ sky130_fd_sc_hd__or2b_1
XFILLER_0_138_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__14212__A2 _02138_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13421_ _05950_ VGND VGND VPWR VPWR _05951_ sky130_fd_sc_hd__inv_2
X_10633_ _02896_ _02897_ _02900_ VGND VGND VPWR VPWR _02902_ sky130_fd_sc_hd__nor3_1
XANTENNA__12223__A1 _00778_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12223__B2 _00783_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13352_ _05341_ _05347_ _05874_ VGND VGND VPWR VPWR _05875_ sky130_fd_sc_hd__and3_1
XFILLER_0_106_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10564_ _00818_ _02758_ _02818_ _02825_ VGND VGND VPWR VPWR _02826_ sky130_fd_sc_hd__a31o_1
XFILLER_0_106_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12303_ _01288_ _02187_ _02189_ _00416_ VGND VGND VPWR VPWR _04738_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_106_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13283_ _05786_ _05802_ _05805_ VGND VGND VPWR VPWR _05806_ sky130_fd_sc_hd__a21oi_1
X_10495_ _00636_ _02735_ _02731_ _00526_ VGND VGND VPWR VPWR _02750_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12234_ _00778_ _01178_ _01248_ _00783_ VGND VGND VPWR VPWR _04662_ sky130_fd_sc_hd__a22o_1
XANTENNA__08699__B _00784_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12165_ _04575_ _04580_ _04585_ _04553_ VGND VGND VPWR VPWR _04586_ sky130_fd_sc_hd__o211a_1
X_11116_ _03431_ _02581_ _03432_ VGND VGND VPWR VPWR _03434_ sky130_fd_sc_hd__a21o_1
X_12096_ _04508_ _04509_ VGND VGND VPWR VPWR _04511_ sky130_fd_sc_hd__nor2_2
XFILLER_0_127_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07108__B _00300_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11047_ _02574_ _03357_ VGND VGND VPWR VPWR _03358_ sky130_fd_sc_hd__nor2_1
Xinput9 a[17] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__buf_4
XANTENNA__09604__A _06417_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_524 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12998_ _05475_ _05484_ VGND VGND VPWR VPWR _05503_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07124__A net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11949_ _04346_ _04348_ VGND VGND VPWR VPWR _04349_ sky130_fd_sc_hd__or2_1
XFILLER_0_143_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08130__A2 _07075_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13619_ _06133_ _06167_ VGND VGND VPWR VPWR _06168_ sky130_fd_sc_hd__and2_1
XANTENNA__12214__A1 _01507_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13499__C _03687_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12214__B2 _00605_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07140_ net59 VGND VGND VPWR VPWR _00901_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_82_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10776__B2 _02116_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12205__A _00374_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07973_ _07008_ _07016_ VGND VGND VPWR VPWR _00017_ sky130_fd_sc_hd__and2_1
XANTENNA__09146__A1 _01295_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09712_ _02160_ _06461_ _01508_ _01504_ VGND VGND VPWR VPWR _01893_ sky130_fd_sc_hd__and4_1
XANTENNA__09146__B2 _01405_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09643_ _01255_ _01571_ _01817_ VGND VGND VPWR VPWR _01818_ sky130_fd_sc_hd__nor3_1
XFILLER_0_96_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09574_ _01740_ _01741_ VGND VGND VPWR VPWR _01742_ sky130_fd_sc_hd__xnor2_1
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08525_ _00579_ _00593_ VGND VGND VPWR VPWR _00594_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08456_ _00516_ _00518_ VGND VGND VPWR VPWR _00520_ sky130_fd_sc_hd__nor2_1
XFILLER_0_65_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07407_ _03784_ _03817_ VGND VGND VPWR VPWR _03828_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_135_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08387_ _04081_ _00373_ _04213_ _04202_ VGND VGND VPWR VPWR _00444_ sky130_fd_sc_hd__a31o_1
XANTENNA__07880__A1 _00891_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07338_ _03059_ VGND VGND VPWR VPWR _03070_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_60_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_755 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11003__B _04598_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07269_ _02291_ _02302_ VGND VGND VPWR VPWR _02313_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_835 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09008_ _03004_ _00113_ _00114_ _00095_ VGND VGND VPWR VPWR _01123_ sky130_fd_sc_hd__a22oi_2
X_10280_ _02513_ _02514_ VGND VGND VPWR VPWR _02515_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11192__A1 _01156_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13970_ _06537_ _06540_ VGND VGND VPWR VPWR _06554_ sky130_fd_sc_hd__nand2_1
X_12921_ _05416_ _05319_ _05312_ VGND VGND VPWR VPWR _05418_ sky130_fd_sc_hd__and3_1
XTAP_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12852_ _01586_ _02306_ _02305_ _00574_ VGND VGND VPWR VPWR _05342_ sky130_fd_sc_hd__a22oi_2
XANTENNA__11392__C _01179_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11803_ _04186_ _02677_ _04187_ VGND VGND VPWR VPWR _04188_ sky130_fd_sc_hd__and3_1
XFILLER_0_139_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12783_ _05264_ _05265_ VGND VGND VPWR VPWR _05266_ sky130_fd_sc_hd__xor2_1
XTAP_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12995__A2 _02008_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11734_ _02630_ _04111_ VGND VGND VPWR VPWR _04112_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_139_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09860__A2 _02039_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11665_ _06885_ _01601_ VGND VGND VPWR VPWR _04036_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_763 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13404_ _03414_ _01956_ _03687_ _04714_ VGND VGND VPWR VPWR _05932_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10616_ _01472_ _01060_ _02882_ _02867_ VGND VGND VPWR VPWR _02884_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_36_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11596_ _03776_ _03959_ VGND VGND VPWR VPWR _03961_ sky130_fd_sc_hd__or2_1
XFILLER_0_52_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13335_ _00745_ _02724_ _02728_ _00914_ VGND VGND VPWR VPWR _05856_ sky130_fd_sc_hd__a22o_1
XANTENNA__07623__A1 _02007_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10547_ _00819_ _00818_ _02725_ _02730_ VGND VGND VPWR VPWR _02808_ sky130_fd_sc_hd__nand4_1
XFILLER_0_122_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13266_ _05760_ _05788_ _05789_ VGND VGND VPWR VPWR _05791_ sky130_fd_sc_hd__a21o_1
XFILLER_0_51_298 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10478_ _01472_ _02726_ _02731_ _00636_ VGND VGND VPWR VPWR _02732_ sky130_fd_sc_hd__a22o_1
XANTENNA__08179__A2 _00219_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12217_ _00458_ _03750_ _04643_ _04639_ VGND VGND VPWR VPWR _04644_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_110_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13197_ _05199_ _05721_ VGND VGND VPWR VPWR _05722_ sky130_fd_sc_hd__xnor2_2
XANTENNA__11567__C _01179_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12148_ _04558_ _04559_ _04561_ VGND VGND VPWR VPWR _04568_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07119__A _00661_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12079_ _03984_ _04404_ VGND VGND VPWR VPWR _04492_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_79_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08351__A2 _00381_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08892__B _00144_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08310_ _00233_ _00239_ _00359_ _00244_ VGND VGND VPWR VPWR _00360_ sky130_fd_sc_hd__o211ai_4
XANTENNA__07789__A net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09290_ _01428_ _01431_ VGND VGND VPWR VPWR _01432_ sky130_fd_sc_hd__xnor2_4
XANTENNA__12986__A2 _05487_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08241_ _00283_ _00284_ VGND VGND VPWR VPWR _00285_ sky130_fd_sc_hd__and2_1
XFILLER_0_144_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08172_ _00208_ _00215_ VGND VGND VPWR VPWR _00216_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_27_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09603__A2 _00415_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07123_ net55 VGND VGND VPWR VPWR _00716_ sky130_fd_sc_hd__buf_6
XFILLER_0_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput110 net110 VGND VGND VPWR VPWR prod[50] sky130_fd_sc_hd__clkbuf_4
XANTENNA__08413__A _02149_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07955__C _00388_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput121 net121 VGND VGND VPWR VPWR prod[60] sky130_fd_sc_hd__buf_6
XFILLER_0_63_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12580__D _02304_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08132__B _00175_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09119__A1 _00344_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07956_ _07084_ VGND VGND VPWR VPWR _00000_ sky130_fd_sc_hd__inv_2
X_07887_ _07009_ _07015_ VGND VGND VPWR VPWR _07016_ sky130_fd_sc_hd__xor2_1
X_09626_ _01797_ _01607_ _01798_ VGND VGND VPWR VPWR _01800_ sky130_fd_sc_hd__a21o_1
XFILLER_0_97_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09557_ _00843_ _00844_ _00635_ _07040_ VGND VGND VPWR VPWR _01724_ sky130_fd_sc_hd__and4_1
XFILLER_0_38_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08508_ _02138_ _00415_ _00575_ _00333_ VGND VGND VPWR VPWR _00576_ sky130_fd_sc_hd__a22o_1
X_09488_ _01434_ _00898_ _01433_ _01636_ VGND VGND VPWR VPWR _01648_ sky130_fd_sc_hd__or4bb_4
XFILLER_0_38_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08439_ _00499_ _00500_ VGND VGND VPWR VPWR _00501_ sky130_fd_sc_hd__nor2_1
XFILLER_0_135_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_828 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11450_ _03797_ _03799_ _03794_ VGND VGND VPWR VPWR _03800_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_92_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10401_ _05445_ _05467_ _01246_ VGND VGND VPWR VPWR _02648_ sky130_fd_sc_hd__and3_1
XFILLER_0_116_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11381_ _01312_ _03699_ _03703_ _03702_ VGND VGND VPWR VPWR _03724_ sky130_fd_sc_hd__a31o_1
XFILLER_0_21_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13120_ _05634_ _05636_ VGND VGND VPWR VPWR _05637_ sky130_fd_sc_hd__nor2_1
X_10332_ _02570_ _02571_ VGND VGND VPWR VPWR _02572_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08323__A _00373_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13051_ _05557_ _05560_ VGND VGND VPWR VPWR _05561_ sky130_fd_sc_hd__nand2_2
X_10263_ _02251_ _02284_ _02288_ _02292_ VGND VGND VPWR VPWR _02496_ sky130_fd_sc_hd__and4bb_2
XANTENNA__07584__D _02664_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12002_ _04357_ _04385_ _04386_ _04387_ VGND VGND VPWR VPWR _04407_ sky130_fd_sc_hd__and4_1
X_10194_ _02410_ _02420_ VGND VGND VPWR VPWR _02421_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_17_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13953_ _06221_ _06534_ VGND VGND VPWR VPWR _06535_ sky130_fd_sc_hd__xnor2_1
X_12904_ _05397_ _05398_ VGND VGND VPWR VPWR _05399_ sky130_fd_sc_hd__and2_1
X_13884_ _06392_ _06458_ VGND VGND VPWR VPWR _06459_ sky130_fd_sc_hd__or2_1
XFILLER_0_69_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12835_ _00916_ _01933_ _05282_ VGND VGND VPWR VPWR _05323_ sky130_fd_sc_hd__and3_1
XTAP_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08097__A1 _04917_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12766_ _05245_ _04654_ _04659_ _05246_ VGND VGND VPWR VPWR _05248_ sky130_fd_sc_hd__nand4_2
XTAP_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09833__A2 _00390_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07402__A _03762_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11717_ _04075_ _04080_ VGND VGND VPWR VPWR _04094_ sky130_fd_sc_hd__nor2_1
X_12697_ _05161_ _05165_ VGND VGND VPWR VPWR _05172_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_126_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_839 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11648_ _03728_ _04017_ VGND VGND VPWR VPWR _04018_ sky130_fd_sc_hd__xor2_1
XFILLER_0_114_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput12 a[1] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__buf_12
XFILLER_0_141_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput23 a[2] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__buf_8
Xinput34 b[10] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__buf_4
XFILLER_0_142_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput45 b[20] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__buf_4
X_11579_ _03909_ _03939_ _03907_ VGND VGND VPWR VPWR _03942_ sky130_fd_sc_hd__a21bo_1
Xinput56 b[30] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09329__A _00544_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13318_ _05839_ VGND VGND VPWR VPWR _05840_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13249_ _02713_ _05579_ _05768_ VGND VGND VPWR VPWR _05775_ sky130_fd_sc_hd__nand3_1
XFILLER_0_20_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07810_ _06527_ _06648_ _06936_ _06938_ VGND VGND VPWR VPWR _06939_ sky130_fd_sc_hd__a211o_1
X_08790_ _00877_ _00884_ VGND VGND VPWR VPWR _00885_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07741_ _06755_ _06869_ VGND VGND VPWR VPWR _06870_ sky130_fd_sc_hd__nand2_1
XANTENNA__09064__A _00344_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07672_ _06712_ net179 VGND VGND VPWR VPWR _06723_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09411_ net19 VGND VGND VPWR VPWR _01564_ sky130_fd_sc_hd__buf_2
XANTENNA__12408__A1 _04059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09342_ _01444_ VGND VGND VPWR VPWR _01488_ sky130_fd_sc_hd__inv_2
XANTENNA__10419__B1 _02133_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09273_ _01412_ VGND VGND VPWR VPWR _01413_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__11631__A2 _01957_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_817 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08224_ _00101_ VGND VGND VPWR VPWR _00268_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_74_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09588__A1 _00991_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_226 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08155_ _00196_ _00198_ VGND VGND VPWR VPWR _00199_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10673__A _00293_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13687__C _02725_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07106_ _00519_ VGND VGND VPWR VPWR _00530_ sky130_fd_sc_hd__buf_4
X_08086_ _00128_ _00129_ VGND VGND VPWR VPWR _00130_ sky130_fd_sc_hd__nor2_1
XANTENNA__08260__A1 _00138_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08260__B2 _06417_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08988_ _01099_ _01100_ VGND VGND VPWR VPWR _01101_ sky130_fd_sc_hd__nand2_1
X_07939_ _06909_ _07067_ VGND VGND VPWR VPWR _07068_ sky130_fd_sc_hd__xnor2_1
X_10950_ _00143_ _04906_ _01508_ _01504_ VGND VGND VPWR VPWR _03251_ sky130_fd_sc_hd__and4_1
XANTENNA__07523__B1 _02960_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09609_ _02040_ _01600_ _01598_ _01597_ _00415_ VGND VGND VPWR VPWR _01781_ sky130_fd_sc_hd__a32o_1
X_10881_ _03082_ _03091_ VGND VGND VPWR VPWR _03175_ sky130_fd_sc_hd__and2_1
XFILLER_0_85_419 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08963__D net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09421__B _00742_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12620_ _01289_ _01061_ _01414_ _01188_ VGND VGND VPWR VPWR _05087_ sky130_fd_sc_hd__a22oi_1
XANTENNA__09276__B1 _01415_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11670__C _03718_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08318__A _00354_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12485__D _00741_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12551_ _00376_ _01188_ _01289_ _00380_ VGND VGND VPWR VPWR _05011_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_108_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11622__A2 _01957_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11502_ _03855_ _03856_ VGND VGND VPWR VPWR _03857_ sky130_fd_sc_hd__or2b_1
XFILLER_0_109_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12482_ _00777_ _03729_ _03762_ _00612_ VGND VGND VPWR VPWR _04935_ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12782__B _01412_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11433_ _03747_ _03756_ VGND VGND VPWR VPWR _03781_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_123_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14221_ _00405_ _06805_ VGND VGND VPWR VPWR _06806_ sky130_fd_sc_hd__nand2_1
XANTENNA__07876__B _07004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14152_ _06726_ _06749_ VGND VGND VPWR VPWR _06751_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11364_ _01312_ _03680_ VGND VGND VPWR VPWR _03705_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13103_ _04032_ VGND VGND VPWR VPWR _05618_ sky130_fd_sc_hd__inv_2
XFILLER_0_132_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10315_ _05192_ net45 _02356_ _02224_ _01506_ VGND VGND VPWR VPWR _02553_ sky130_fd_sc_hd__a32o_1
XFILLER_0_104_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14083_ _06102_ _06650_ _06676_ VGND VGND VPWR VPWR _06677_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_131_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11295_ _02862_ _02908_ _02859_ VGND VGND VPWR VPWR _03630_ sky130_fd_sc_hd__a21bo_1
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13034_ _05532_ _05539_ _05541_ VGND VGND VPWR VPWR _05542_ sky130_fd_sc_hd__a21o_1
X_10246_ _02476_ _02477_ VGND VGND VPWR VPWR _02479_ sky130_fd_sc_hd__or2_1
XANTENNA__09200__B1 _00298_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10177_ _00101_ _06733_ _03685_ _00423_ VGND VGND VPWR VPWR _02403_ sky130_fd_sc_hd__and4_1
XANTENNA__12022__B _06450_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13936_ _06499_ _06515_ VGND VGND VPWR VPWR _06517_ sky130_fd_sc_hd__nand2_1
XANTENNA__07514__B1 net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13867_ _06429_ _06440_ VGND VGND VPWR VPWR _06441_ sky130_fd_sc_hd__and2_1
XFILLER_0_147_819 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12818_ _05260_ _05261_ _05262_ _05303_ VGND VGND VPWR VPWR _05305_ sky130_fd_sc_hd__o31ai_2
XFILLER_0_146_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13798_ _02188_ _02190_ _03684_ _03680_ VGND VGND VPWR VPWR _06365_ sky130_fd_sc_hd__and4_1
XANTENNA__08228__A _06461_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12395__D _00571_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12749_ _05224_ _05228_ VGND VGND VPWR VPWR _05229_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_56_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10821__B1 net57 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09985__C _02187_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_861 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07786__B _04378_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10493__A _02247_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_719 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09059__A _01178_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09960_ _02163_ _02164_ VGND VGND VPWR VPWR _02165_ sky130_fd_sc_hd__and2b_1
XFILLER_0_122_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08911_ _01013_ _01016_ VGND VGND VPWR VPWR _01017_ sky130_fd_sc_hd__xnor2_1
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09891_ _03070_ _02088_ _01983_ _01984_ VGND VGND VPWR VPWR _02089_ sky130_fd_sc_hd__a31o_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08842_ _00729_ _00763_ VGND VGND VPWR VPWR _00941_ sky130_fd_sc_hd__nand2_1
XANTENNA__12213__A _00605_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07307__A _01470_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08773_ _00864_ _00865_ VGND VGND VPWR VPWR _00866_ sky130_fd_sc_hd__nor2_2
XFILLER_0_109_82 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07724_ _02259_ _03543_ _00508_ _02171_ VGND VGND VPWR VPWR _06853_ sky130_fd_sc_hd__a22oi_1
XANTENNA__10104__A2 _01410_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07655_ _06505_ _06516_ _06197_ _06230_ VGND VGND VPWR VPWR _06538_ sky130_fd_sc_hd__a211oi_1
XANTENNA__10668__A _02982_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12586__C _02158_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07586_ _02029_ _05588_ _05753_ _05780_ VGND VGND VPWR VPWR _05790_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_48_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09325_ _00654_ _00635_ _07040_ _00844_ VGND VGND VPWR VPWR _01469_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09256_ _01380_ _01393_ VGND VGND VPWR VPWR _01395_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_106_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08207_ _07083_ _00183_ _00189_ _00249_ _00250_ VGND VGND VPWR VPWR _00251_ sky130_fd_sc_hd__a221o_2
XFILLER_0_7_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09187_ _01123_ _01126_ _01124_ VGND VGND VPWR VPWR _01319_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_90_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08138_ _00180_ _00181_ VGND VGND VPWR VPWR _00182_ sky130_fd_sc_hd__and2b_1
XFILLER_0_43_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10553__D _02723_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11011__B _00604_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08069_ _00112_ VGND VGND VPWR VPWR _00113_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_113_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10100_ _01933_ _02172_ _02317_ VGND VGND VPWR VPWR _02318_ sky130_fd_sc_hd__and3_1
X_11080_ _03391_ _03393_ VGND VGND VPWR VPWR _03394_ sky130_fd_sc_hd__nand2_1
X_10031_ _01753_ VGND VGND VPWR VPWR _02243_ sky130_fd_sc_hd__inv_2
XANTENNA__09416__B _01564_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07217__A _00672_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09135__C _03773_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11982_ _04382_ _04383_ _04384_ VGND VGND VPWR VPWR _04385_ sky130_fd_sc_hd__nand3_2
XFILLER_0_98_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09432__A _00159_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13721_ _06259_ _06279_ VGND VGND VPWR VPWR _06280_ sky130_fd_sc_hd__and2_1
X_10933_ _03223_ _03231_ VGND VGND VPWR VPWR _03232_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13652_ _06195_ VGND VGND VPWR VPWR _06204_ sky130_fd_sc_hd__inv_2
X_10864_ _02528_ _02531_ _03155_ VGND VGND VPWR VPWR _03156_ sky130_fd_sc_hd__a21o_1
XFILLER_0_85_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12603_ _05066_ _05067_ VGND VGND VPWR VPWR _05068_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_94_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13583_ _03785_ _02858_ _03783_ _02856_ VGND VGND VPWR VPWR _06128_ sky130_fd_sc_hd__a22o_1
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10795_ _02259_ _02171_ _02758_ _02169_ VGND VGND VPWR VPWR _03080_ sky130_fd_sc_hd__and4_1
XFILLER_0_54_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12534_ _04989_ _04988_ VGND VGND VPWR VPWR _04992_ sky130_fd_sc_hd__nor2_1
XFILLER_0_109_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13348__A2 _02306_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12465_ _04860_ _04868_ VGND VGND VPWR VPWR _04916_ sky130_fd_sc_hd__and2_1
XANTENNA__11359__A1 _01155_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_680 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14204_ _02324_ VGND VGND VPWR VPWR _06795_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11416_ _03760_ _03761_ _03758_ VGND VGND VPWR VPWR _03763_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_1_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12396_ _00374_ _01272_ _04838_ _04839_ VGND VGND VPWR VPWR _04841_ sky130_fd_sc_hd__a31o_1
XFILLER_0_50_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14135_ _02743_ _04014_ _02742_ _04013_ VGND VGND VPWR VPWR _06732_ sky130_fd_sc_hd__nand4_1
X_11347_ _03686_ VGND VGND VPWR VPWR _03687_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14066_ _06099_ _06656_ VGND VGND VPWR VPWR _06659_ sky130_fd_sc_hd__or2_1
X_11278_ _03602_ _03611_ VGND VGND VPWR VPWR _03612_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13017_ _05519_ _05523_ VGND VGND VPWR VPWR _05524_ sky130_fd_sc_hd__xor2_4
X_10229_ _01394_ net21 net22 _01470_ VGND VGND VPWR VPWR _02460_ sky130_fd_sc_hd__a22o_1
XANTENNA__07127__A _00541_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13919_ _06486_ _06497_ VGND VGND VPWR VPWR _06498_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10488__A _02736_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07440_ net43 VGND VGND VPWR VPWR _04191_ sky130_fd_sc_hd__buf_4
XFILLER_0_9_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07371_ _03114_ _03422_ VGND VGND VPWR VPWR _03433_ sky130_fd_sc_hd__xnor2_2
XANTENNA__13799__A _02187_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09110_ _00984_ _01048_ VGND VGND VPWR VPWR _01235_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09041_ _01157_ _01158_ VGND VGND VPWR VPWR _01159_ sky130_fd_sc_hd__nand2_2
XFILLER_0_26_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12853__D _02305_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap142 _03701_ VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09943_ _02006_ _02028_ _01980_ VGND VGND VPWR VPWR _02146_ sky130_fd_sc_hd__a21o_1
XFILLER_0_111_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10670__B _00151_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13039__A _05541_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13511__A2 _02722_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09874_ _02068_ _02069_ VGND VGND VPWR VPWR _02070_ sky130_fd_sc_hd__or2b_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08825_ _01996_ _03762_ VGND VGND VPWR VPWR _00922_ sky130_fd_sc_hd__nand2_1
XANTENNA__13981__B _06552_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12878__A _01507_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08756_ _00669_ _00674_ _00846_ VGND VGND VPWR VPWR _00848_ sky130_fd_sc_hd__and3_1
XTAP_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07707_ _06834_ _06835_ VGND VGND VPWR VPWR _06836_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_68_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08687_ _00769_ _00771_ VGND VGND VPWR VPWR _00772_ sky130_fd_sc_hd__xnor2_1
XTAP_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07638_ _05654_ _06329_ VGND VGND VPWR VPWR _06351_ sky130_fd_sc_hd__and2_1
XTAP_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_430 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13578__A2 _02858_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07569_ _01361_ _05566_ _05599_ VGND VGND VPWR VPWR _05610_ sky130_fd_sc_hd__and3_1
XFILLER_0_119_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11589__A1 _01155_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_411 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09308_ _00844_ _00819_ VGND VGND VPWR VPWR _01451_ sky130_fd_sc_hd__nand2_1
XANTENNA__07257__A2 _02138_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10580_ _00143_ _02306_ _02305_ _04906_ VGND VGND VPWR VPWR _02844_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07500__A net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09239_ _01072_ _01078_ _01374_ VGND VGND VPWR VPWR _01376_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_51_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12250_ _00375_ _03738_ VGND VGND VPWR VPWR _04680_ sky130_fd_sc_hd__nand2_1
XFILLER_0_121_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10013__A1 _03015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11201_ _03524_ _03526_ VGND VGND VPWR VPWR _03527_ sky130_fd_sc_hd__xnor2_4
XANTENNA__10013__B2 _00388_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11957__A _06417_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12181_ _03548_ _03549_ VGND VGND VPWR VPWR _04604_ sky130_fd_sc_hd__and2_1
XANTENNA__10564__A2 _02758_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11132_ _03049_ _03016_ _03045_ VGND VGND VPWR VPWR _03451_ sky130_fd_sc_hd__or3_1
XANTENNA__11676__B _00268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11063_ _03333_ _03374_ VGND VGND VPWR VPWR _03375_ sky130_fd_sc_hd__nor2_1
XANTENNA__11395__C _06765_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10014_ _00366_ _02971_ net46 VGND VGND VPWR VPWR _02224_ sky130_fd_sc_hd__and3_1
XANTENNA__09182__A2 _00636_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09162__A _03070_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11965_ _04292_ _04294_ _04364_ VGND VGND VPWR VPWR _04366_ sky130_fd_sc_hd__nor3_1
XANTENNA_output116_A net116 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12300__B _02426_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13704_ _06250_ _06260_ VGND VGND VPWR VPWR _06261_ sky130_fd_sc_hd__nor2_1
X_10916_ _03194_ _03196_ VGND VGND VPWR VPWR _03214_ sky130_fd_sc_hd__xnor2_1
X_11896_ _04148_ _04149_ VGND VGND VPWR VPWR _04291_ sky130_fd_sc_hd__and2b_1
XFILLER_0_67_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13635_ _06180_ _06184_ VGND VGND VPWR VPWR _06185_ sky130_fd_sc_hd__and2b_1
XFILLER_0_132_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10847_ _03116_ _03118_ _03137_ _03112_ VGND VGND VPWR VPWR _03138_ sky130_fd_sc_hd__a211o_1
XFILLER_0_67_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13566_ _06108_ _06079_ VGND VGND VPWR VPWR _06110_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_137_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10778_ _06937_ _02169_ _03060_ _03061_ VGND VGND VPWR VPWR _03062_ sky130_fd_sc_hd__a31o_1
XFILLER_0_82_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08506__A _00572_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08996__A2 _01108_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12517_ _04962_ _04964_ VGND VGND VPWR VPWR _04974_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_124_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13497_ _06009_ _03684_ VGND VGND VPWR VPWR _06034_ sky130_fd_sc_hd__nand2_1
XANTENNA__08225__B _02149_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12448_ _04889_ _04897_ VGND VGND VPWR VPWR _04898_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_112_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10004__A1 _04598_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10004__B2 _05192_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12379_ _04794_ _04797_ VGND VGND VPWR VPWR _04822_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14118_ _06654_ _06713_ VGND VGND VPWR VPWR _06715_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_560 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07783__C _00355_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10490__B _02742_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14049_ _06638_ _06640_ VGND VGND VPWR VPWR _06641_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_5_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08610_ _00316_ _00510_ _00509_ VGND VGND VPWR VPWR _00688_ sky130_fd_sc_hd__o21ba_1
X_09590_ _01754_ _01758_ _01718_ VGND VGND VPWR VPWR _01760_ sky130_fd_sc_hd__a21oi_2
X_08541_ _04103_ VGND VGND VPWR VPWR _00612_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_49_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_50 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08472_ _00531_ _00536_ VGND VGND VPWR VPWR _00537_ sky130_fd_sc_hd__xor2_1
XANTENNA__08684__A1 _00639_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08684__B2 _00563_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07423_ _03982_ _03993_ VGND VGND VPWR VPWR _04004_ sky130_fd_sc_hd__or2b_4
XFILLER_0_92_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07354_ _03224_ net147 VGND VGND VPWR VPWR _03246_ sky130_fd_sc_hd__xor2_2
XANTENNA__08416__A _06483_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07285_ _00847_ _01864_ VGND VGND VPWR VPWR _02489_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08135__B _00002_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11991__A1 _00530_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09024_ _03543_ _00298_ _01138_ VGND VGND VPWR VPWR _01140_ sky130_fd_sc_hd__and3_1
XFILLER_0_103_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12880__B _02120_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10546__A2 _02169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09247__A _02664_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07411__A2 _03685_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07693__C _06819_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09926_ _01818_ _01973_ _01972_ VGND VGND VPWR VPWR _02128_ sky130_fd_sc_hd__a21o_1
XANTENNA__13496__A1 _01415_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09857_ _01760_ _02041_ _02042_ VGND VGND VPWR VPWR _02052_ sky130_fd_sc_hd__and3b_2
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08808_ _02127_ _00734_ VGND VGND VPWR VPWR _00904_ sky130_fd_sc_hd__nand2_1
X_09788_ _02456_ _01180_ _01976_ VGND VGND VPWR VPWR _01977_ sky130_fd_sc_hd__and3_1
XTAP_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08739_ _00827_ _00828_ VGND VGND VPWR VPWR _00829_ sky130_fd_sc_hd__xor2_1
XTAP_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07478__A2 net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ _04113_ _04129_ VGND VGND VPWR VPWR _04130_ sky130_fd_sc_hd__nor2_1
XTAP_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10701_ _00095_ _01059_ VGND VGND VPWR VPWR _02977_ sky130_fd_sc_hd__nand2_1
XTAP_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10856__A _06483_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11681_ _04047_ _04053_ VGND VGND VPWR VPWR _04054_ sky130_fd_sc_hd__xor2_1
XTAP_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13420_ _01061_ _01181_ _01414_ _01250_ VGND VGND VPWR VPWR _05950_ sky130_fd_sc_hd__and4_1
X_10632_ _02896_ _02897_ _02900_ VGND VGND VPWR VPWR _02901_ sky130_fd_sc_hd__o21a_1
XANTENNA__12223__A2 _01248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08326__A _04059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_403 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10563_ _02824_ VGND VGND VPWR VPWR _02825_ sky130_fd_sc_hd__inv_2
X_13351_ _05870_ _05873_ VGND VGND VPWR VPWR _05874_ sky130_fd_sc_hd__xor2_1
XFILLER_0_106_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12302_ _00415_ _00575_ _01664_ _01505_ VGND VGND VPWR VPWR _04737_ sky130_fd_sc_hd__and4_1
XFILLER_0_106_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13282_ _05797_ _05801_ _05804_ VGND VGND VPWR VPWR _05805_ sky130_fd_sc_hd__a21o_1
X_10494_ _02747_ _02748_ VGND VGND VPWR VPWR _02749_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_32_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12233_ _04659_ _04660_ VGND VGND VPWR VPWR _04661_ sky130_fd_sc_hd__nand2_1
XANTENNA__10591__A _02855_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12164_ _04581_ _04584_ _04403_ _04454_ VGND VGND VPWR VPWR _04585_ sky130_fd_sc_hd__and4_1
XFILLER_0_20_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08061__A _05588_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11115_ _02545_ _02578_ VGND VGND VPWR VPWR _03432_ sky130_fd_sc_hd__and2b_1
X_12095_ _04507_ _04436_ _04439_ VGND VGND VPWR VPWR _04509_ sky130_fd_sc_hd__nor3_1
X_11046_ _03353_ _03354_ VGND VGND VPWR VPWR _03357_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09604__B _00138_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12997_ _05493_ _05494_ _05495_ _05501_ VGND VGND VPWR VPWR _05502_ sky130_fd_sc_hd__a31o_1
XFILLER_0_143_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11948_ _04347_ _04344_ VGND VGND VPWR VPWR _04348_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11879_ _04091_ _04100_ VGND VGND VPWR VPWR _04272_ sky130_fd_sc_hd__nand2_1
XANTENNA__12684__C _05150_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13618_ _06140_ _06143_ _06166_ VGND VGND VPWR VPWR _06167_ sky130_fd_sc_hd__a21o_1
XANTENNA__08418__A1 _06472_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12214__A2 _01179_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07140__A net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13549_ _06089_ _06090_ VGND VGND VPWR VPWR _06091_ sky130_fd_sc_hd__nor2_1
XANTENNA__10776__A2 _02723_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09067__A _00416_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12205__B _00784_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07972_ _00014_ _00015_ VGND VGND VPWR VPWR _00016_ sky130_fd_sc_hd__or2_1
X_09711_ _06461_ _01508_ _01505_ _02160_ VGND VGND VPWR VPWR _01892_ sky130_fd_sc_hd__a22o_1
XANTENNA__09146__A2 _01272_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09642_ _01813_ _01816_ VGND VGND VPWR VPWR _01817_ sky130_fd_sc_hd__xnor2_1
X_09573_ _01457_ _01458_ _01462_ _01334_ VGND VGND VPWR VPWR _01741_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_78_834 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08524_ _00589_ _00592_ VGND VGND VPWR VPWR _00593_ sky130_fd_sc_hd__xor2_1
XFILLER_0_77_355 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08455_ _00291_ _00302_ _00517_ VGND VGND VPWR VPWR _00518_ sky130_fd_sc_hd__a21o_1
XFILLER_0_93_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07406_ _03795_ _03806_ VGND VGND VPWR VPWR _03817_ sky130_fd_sc_hd__and2b_1
X_08386_ _04246_ _04290_ VGND VGND VPWR VPWR _00443_ sky130_fd_sc_hd__nand2_1
XFILLER_0_147_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07880__A2 net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07337_ _02018_ VGND VGND VPWR VPWR _03059_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__11413__B1 _01248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12891__A _00779_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07268_ net156 _01700_ _01788_ VGND VGND VPWR VPWR _02302_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11003__C _01368_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_847 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09007_ _01008_ _01010_ VGND VGND VPWR VPWR _01122_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07199_ _01273_ _01317_ _01262_ VGND VGND VPWR VPWR _01547_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_131_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11192__A2 _01108_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09909_ _02086_ _02108_ VGND VGND VPWR VPWR _02109_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13227__A _05424_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12920_ _05319_ _05312_ _05416_ VGND VGND VPWR VPWR _05417_ sky130_fd_sc_hd__a21oi_4
XTAP_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12851_ _02857_ _05091_ _05264_ _05265_ VGND VGND VPWR VPWR _05341_ sky130_fd_sc_hd__o2bb2ai_1
XTAP_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11392__D _01254_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11802_ _04172_ _04177_ VGND VGND VPWR VPWR _04187_ sky130_fd_sc_hd__xnor2_1
XTAP_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_130 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12782_ _01600_ _01412_ VGND VGND VPWR VPWR _05265_ sky130_fd_sc_hd__nand2_1
XTAP_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11733_ _04110_ _04078_ VGND VGND VPWR VPWR _04111_ sky130_fd_sc_hd__nor2_1
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10586__A _04895_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11664_ _00575_ _04033_ _04034_ VGND VGND VPWR VPWR _04035_ sky130_fd_sc_hd__a21bo_1
X_13403_ _05929_ _05930_ VGND VGND VPWR VPWR _05931_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10615_ _02866_ VGND VGND VPWR VPWR _02882_ sky130_fd_sc_hd__inv_2
X_11595_ _03774_ _03775_ VGND VGND VPWR VPWR _03959_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13334_ _05327_ _05330_ _05328_ VGND VGND VPWR VPWR _05855_ sky130_fd_sc_hd__o21ba_1
XANTENNA__07623__A2 _05588_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10546_ _00818_ _02169_ _02798_ _02797_ VGND VGND VPWR VPWR _02807_ sky130_fd_sc_hd__a31o_1
XFILLER_0_134_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13265_ _05507_ _05524_ _05593_ _05597_ VGND VGND VPWR VPWR _05789_ sky130_fd_sc_hd__a31o_1
X_10477_ _02730_ VGND VGND VPWR VPWR _02731_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__12306__A _01400_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12216_ _01664_ _01180_ _01249_ _00607_ VGND VGND VPWR VPWR _04643_ sky130_fd_sc_hd__a22oi_1
X_13196_ _05198_ _05200_ VGND VGND VPWR VPWR _05721_ sky130_fd_sc_hd__nand2_1
XFILLER_0_121_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11567__D _01254_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12147_ _04566_ VGND VGND VPWR VPWR _04567_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12078_ _04403_ _04454_ _04486_ _04490_ VGND VGND VPWR VPWR _04491_ sky130_fd_sc_hd__a31oi_2
X_11029_ _00158_ _04037_ _03336_ _03337_ VGND VGND VPWR VPWR _03338_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10143__B1 _00782_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_300 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11880__A _00257_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_826 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10496__A _00636_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08240_ _00128_ _00131_ VGND VGND VPWR VPWR _00284_ sky130_fd_sc_hd__or2b_1
XFILLER_0_28_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08171_ _00210_ _00214_ VGND VGND VPWR VPWR _00215_ sky130_fd_sc_hd__xnor2_1
X_07122_ net58 VGND VGND VPWR VPWR _00705_ sky130_fd_sc_hd__buf_8
XFILLER_0_70_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13600__A _01061_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput100 net100 VGND VGND VPWR VPWR prod[41] sky130_fd_sc_hd__clkbuf_4
Xoutput111 net111 VGND VGND VPWR VPWR prod[51] sky130_fd_sc_hd__clkbuf_4
XANTENNA__07955__D _03004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput122 net122 VGND VGND VPWR VPWR prod[61] sky130_fd_sc_hd__buf_6
XANTENNA__08413__B _05577_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09119__A2 _01182_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07955_ _03532_ _00497_ _00388_ _03004_ VGND VGND VPWR VPWR _07084_ sky130_fd_sc_hd__and4_1
X_07886_ _07013_ _07014_ VGND VGND VPWR VPWR _07015_ sky130_fd_sc_hd__xnor2_1
X_09625_ _01573_ _01595_ VGND VGND VPWR VPWR _01798_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09556_ _01466_ _01478_ VGND VGND VPWR VPWR _01723_ sky130_fd_sc_hd__nand2_1
XANTENNA__09260__A _02116_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08507_ _00574_ VGND VGND VPWR VPWR _00575_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_38_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09487_ _01433_ _01436_ _01636_ _01643_ _01646_ VGND VGND VPWR VPWR _01647_ sky130_fd_sc_hd__a32oi_4
XANTENNA__07302__A1 _02664_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08438_ _05456_ _05478_ _00142_ _04862_ VGND VGND VPWR VPWR _00500_ sky130_fd_sc_hd__and4_1
XFILLER_0_81_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08369_ _03850_ _00423_ net10 _01306_ VGND VGND VPWR VPWR _00424_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_135_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10400_ _02444_ _02446_ VGND VGND VPWR VPWR _02647_ sky130_fd_sc_hd__and2_1
X_11380_ _03711_ _03722_ VGND VGND VPWR VPWR _03723_ sky130_fd_sc_hd__and2b_1
XFILLER_0_21_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10331_ net7 _04048_ VGND VGND VPWR VPWR _02571_ sky130_fd_sc_hd__nand2_1
XANTENNA__11030__A _05027_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13050_ _05549_ _05556_ _05559_ VGND VGND VPWR VPWR _05560_ sky130_fd_sc_hd__o21ai_1
X_10262_ _02491_ _02495_ VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__xor2_1
X_12001_ _04404_ _04405_ VGND VGND VPWR VPWR _04406_ sky130_fd_sc_hd__nor2_1
X_10193_ _02418_ _02419_ VGND VGND VPWR VPWR _02420_ sky130_fd_sc_hd__nand2_1
XFILLER_0_108_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13952_ _06225_ _06224_ VGND VGND VPWR VPWR _06534_ sky130_fd_sc_hd__and2b_1
X_12903_ _05380_ _05396_ VGND VGND VPWR VPWR _05398_ sky130_fd_sc_hd__or2_1
X_13883_ _05935_ _06391_ VGND VGND VPWR VPWR _06458_ sky130_fd_sc_hd__and2_1
XANTENNA__12796__A _00389_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12834_ _05282_ _05283_ VGND VGND VPWR VPWR _05322_ sky130_fd_sc_hd__or2b_1
XTAP_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12765_ _04661_ _04698_ VGND VGND VPWR VPWR _05246_ sky130_fd_sc_hd__or2b_1
XTAP_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13090__A2 _05595_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11716_ _04062_ _04067_ _04074_ VGND VGND VPWR VPWR _04093_ sky130_fd_sc_hd__and3_1
XTAP_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12696_ _05157_ _05158_ _05169_ VGND VGND VPWR VPWR _05171_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_37_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11647_ _02246_ _04013_ _04016_ VGND VGND VPWR VPWR _04017_ sky130_fd_sc_hd__and3_1
XFILLER_0_71_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput13 a[20] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_52_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13420__A _01061_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput24 a[30] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__buf_4
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput35 b[11] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__buf_2
XFILLER_0_107_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput46 b[21] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__buf_4
XFILLER_0_25_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__08514__A _01361_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11578_ _03912_ _03936_ _03940_ VGND VGND VPWR VPWR _03941_ sky130_fd_sc_hd__a21oi_1
Xinput57 b[31] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13317_ _05679_ _05741_ _05747_ VGND VGND VPWR VPWR _05839_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09329__B _01473_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10529_ _02770_ _02785_ _02787_ _02782_ VGND VGND VPWR VPWR _02788_ sky130_fd_sc_hd__o31a_1
X_13248_ _01837_ _02045_ _02274_ _02491_ VGND VGND VPWR VPWR _05774_ sky130_fd_sc_hd__nand4_1
XFILLER_0_122_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12353__A1 _00742_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13179_ _04531_ _04536_ _04490_ VGND VGND VPWR VPWR _05702_ sky130_fd_sc_hd__nand3_1
X_07740_ _06867_ _06868_ VGND VGND VPWR VPWR _06869_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09064__B _01183_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10667__A1 _05192_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07671_ _06680_ _06701_ VGND VGND VPWR VPWR _06712_ sky130_fd_sc_hd__nor2_1
XANTENNA__10667__B2 _02982_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09410_ _01300_ _01301_ _01302_ _01562_ _01256_ VGND VGND VPWR VPWR _01563_ sky130_fd_sc_hd__a32o_2
XFILLER_0_90_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12408__A2 _01272_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10419__A1 _01295_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09341_ _01443_ _01444_ _01486_ VGND VGND VPWR VPWR _01487_ sky130_fd_sc_hd__a21o_1
XANTENNA__10419__B2 _01306_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09272_ _01411_ VGND VGND VPWR VPWR _01412_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_35_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08223_ _00255_ _00266_ VGND VGND VPWR VPWR _00267_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_62_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08154_ _06884_ _00197_ VGND VGND VPWR VPWR _00198_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_132_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10673__B _02855_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13687__D _02728_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07105_ _00508_ VGND VGND VPWR VPWR _00519_ sky130_fd_sc_hd__buf_4
X_08085_ _00032_ _00127_ VGND VGND VPWR VPWR _00129_ sky130_fd_sc_hd__nor2_1
XANTENNA__08260__A2 _04906_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08987_ _01083_ _01097_ VGND VGND VPWR VPWR _01100_ sky130_fd_sc_hd__or2_1
X_07938_ _07065_ _07066_ VGND VGND VPWR VPWR _07067_ sky130_fd_sc_hd__and2b_1
XFILLER_0_97_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07869_ _06986_ _06987_ _06997_ VGND VGND VPWR VPWR _06998_ sky130_fd_sc_hd__a21o_4
XFILLER_0_97_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07523__B2 net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08720__B1 _04873_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09608_ _01585_ VGND VGND VPWR VPWR _01780_ sky130_fd_sc_hd__clkbuf_4
X_10880_ _03172_ _03173_ VGND VGND VPWR VPWR _03174_ sky130_fd_sc_hd__or2_1
XANTENNA__07503__A _01744_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09539_ _00355_ _02960_ net41 _04180_ VGND VGND VPWR VPWR _01704_ sky130_fd_sc_hd__and4_1
XANTENNA__09276__A1 _02051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09276__B2 _00464_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11670__D net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_420 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12550_ _05004_ _05006_ _05009_ VGND VGND VPWR VPWR _05010_ sky130_fd_sc_hd__a21o_1
XFILLER_0_109_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11501_ _03849_ _03852_ VGND VGND VPWR VPWR _03856_ sky130_fd_sc_hd__or2_1
XANTENNA__10830__A1 _04081_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10830__B2 _02727_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12481_ _04820_ _04933_ VGND VGND VPWR VPWR _04934_ sky130_fd_sc_hd__nor2_1
X_14220_ _00404_ VGND VGND VPWR VPWR _06805_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11432_ _03772_ _03778_ _03779_ VGND VGND VPWR VPWR _03780_ sky130_fd_sc_hd__o21a_1
XFILLER_0_80_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14151_ _06726_ _06749_ VGND VGND VPWR VPWR _06750_ sky130_fd_sc_hd__or2_1
X_11363_ _03702_ _03703_ VGND VGND VPWR VPWR _03704_ sky130_fd_sc_hd__and2b_1
XFILLER_0_1_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13102_ _05459_ _05461_ _05462_ _05614_ _05616_ VGND VGND VPWR VPWR _05617_ sky130_fd_sc_hd__o311a_1
X_10314_ _02550_ _02551_ VGND VGND VPWR VPWR _02552_ sky130_fd_sc_hd__xor2_1
X_14082_ _06660_ _06675_ VGND VGND VPWR VPWR _06676_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11294_ _02789_ _03628_ VGND VGND VPWR VPWR _03629_ sky130_fd_sc_hd__nor2_1
XFILLER_0_131_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13033_ _04970_ _04971_ VGND VGND VPWR VPWR _05541_ sky130_fd_sc_hd__xor2_4
XANTENNA__11695__A _06964_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10245_ _02473_ _02475_ VGND VGND VPWR VPWR _02477_ sky130_fd_sc_hd__and2_1
XANTENNA__09200__A1 _00262_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09200__B2 _00263_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10176_ _02400_ VGND VGND VPWR VPWR _02402_ sky130_fd_sc_hd__inv_2
XANTENNA__12022__C _03683_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13935_ _06496_ _06498_ VGND VGND VPWR VPWR _06515_ sky130_fd_sc_hd__or2_1
XANTENNA__07514__A1 net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07514__B2 _00573_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13866_ _05921_ _05926_ _06427_ VGND VGND VPWR VPWR _06440_ sky130_fd_sc_hd__or3_1
XANTENNA__08509__A _01744_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07413__A net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13134__B _05651_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12817_ _05260_ _05261_ _05262_ _05303_ VGND VGND VPWR VPWR _05304_ sky130_fd_sc_hd__or4_4
XFILLER_0_9_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13797_ _06242_ _06253_ _06290_ _06363_ VGND VGND VPWR VPWR _06364_ sky130_fd_sc_hd__nor4_1
XANTENNA__08228__B _00003_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12748_ _05226_ _05227_ VGND VGND VPWR VPWR _05228_ sky130_fd_sc_hd__xnor2_1
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12973__B _05447_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_166 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10821__A1 _00891_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10821__B2 _00989_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10774__A _06494_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12679_ _05136_ _05151_ VGND VGND VPWR VPWR _05152_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09985__D _02189_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12023__B1 _03679_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10493__B _02721_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08910_ _01014_ _01015_ VGND VGND VPWR VPWR _01016_ sky130_fd_sc_hd__xnor2_1
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09890_ _01780_ VGND VGND VPWR VPWR _02088_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_110_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_291 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08841_ _00936_ _00939_ VGND VGND VPWR VPWR _00940_ sky130_fd_sc_hd__xnor2_4
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12213__B _01507_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10014__A _00366_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07307__B _02719_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08772_ _00696_ _00699_ _00863_ VGND VGND VPWR VPWR _00865_ sky130_fd_sc_hd__o21a_1
XANTENNA__13826__A1 _00460_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13826__B2 _01955_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07723_ _02105_ _00650_ _03510_ _00475_ VGND VGND VPWR VPWR _06852_ sky130_fd_sc_hd__and4_1
XFILLER_0_79_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07654_ _06197_ _06230_ _06505_ _06516_ VGND VGND VPWR VPWR _06527_ sky130_fd_sc_hd__o211a_2
XANTENNA__10668__B _05192_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12586__D _02304_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07585_ _05761_ VGND VGND VPWR VPWR _05780_ sky130_fd_sc_hd__inv_2
X_09324_ _00844_ _00654_ _00635_ VGND VGND VPWR VPWR _01468_ sky130_fd_sc_hd__and3_1
XFILLER_0_47_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09255_ _01391_ _01392_ VGND VGND VPWR VPWR _01393_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08206_ _00089_ _00181_ _00180_ VGND VGND VPWR VPWR _00250_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_145_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09186_ _01122_ _01127_ VGND VGND VPWR VPWR _01318_ sky130_fd_sc_hd__or2b_1
XFILLER_0_43_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08137_ _00083_ _00179_ _00178_ VGND VGND VPWR VPWR _00181_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_71_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_411 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08068_ _07010_ VGND VGND VPWR VPWR _00112_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__12317__A1 _00460_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12404__A _00374_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10030_ _02152_ _01948_ _01949_ _02240_ _02241_ VGND VGND VPWR VPWR _02242_ sky130_fd_sc_hd__o41a_2
XANTENNA__09416__C _00311_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09135__D _01260_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11981_ _04232_ _04251_ _04319_ _04288_ VGND VGND VPWR VPWR _04384_ sky130_fd_sc_hd__a211o_1
XANTENNA__10859__A _03268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_556 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13720_ _06247_ _06258_ _06257_ VGND VGND VPWR VPWR _06279_ sky130_fd_sc_hd__o21ai_1
X_10932_ _03225_ _03229_ _03230_ VGND VGND VPWR VPWR _03231_ sky130_fd_sc_hd__o21bai_1
XANTENNA__09432__B _01586_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08329__A _00380_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13651_ _06201_ _06202_ VGND VGND VPWR VPWR _06203_ sky130_fd_sc_hd__or2_1
X_10863_ _05566_ _01058_ _02529_ VGND VGND VPWR VPWR _03155_ sky130_fd_sc_hd__and3_1
XFILLER_0_79_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12602_ _00914_ _01412_ VGND VGND VPWR VPWR _05067_ sky130_fd_sc_hd__nand2_1
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13582_ _06009_ _03785_ _02858_ _03783_ VGND VGND VPWR VPWR _06127_ sky130_fd_sc_hd__nand4_1
XFILLER_0_66_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10794_ _03077_ _03078_ VGND VGND VPWR VPWR _03079_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12533_ _04929_ _04990_ VGND VGND VPWR VPWR _04991_ sky130_fd_sc_hd__xor2_1
XPHY_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10594__A _00145_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12005__B1 _02088_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07680__B1 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12464_ _04821_ _04914_ VGND VGND VPWR VPWR _04915_ sky130_fd_sc_hd__and2_1
X_14203_ _06793_ _06794_ VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__xnor2_4
XFILLER_0_34_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11202__B _03527_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11415_ _06775_ _02119_ VGND VGND VPWR VPWR _03761_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12395_ _00782_ _00613_ _00413_ _00571_ VGND VGND VPWR VPWR _04839_ sky130_fd_sc_hd__and4_1
XFILLER_0_105_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14134_ _04014_ _02742_ _04013_ _02743_ VGND VGND VPWR VPWR _06731_ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11346_ _02135_ VGND VGND VPWR VPWR _03686_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_104_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14065_ _06099_ _06656_ VGND VGND VPWR VPWR _06657_ sky130_fd_sc_hd__nand2_1
X_11277_ _03608_ _03610_ VGND VGND VPWR VPWR _03611_ sky130_fd_sc_hd__and2b_2
XANTENNA__12314__A _00459_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13016_ _05501_ _05521_ VGND VGND VPWR VPWR _05523_ sky130_fd_sc_hd__xnor2_4
X_10228_ net24 VGND VGND VPWR VPWR _02459_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_146_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07127__B _00661_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10159_ _02378_ _02381_ VGND VGND VPWR VPWR _02383_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13918_ _06485_ _06433_ _06482_ VGND VGND VPWR VPWR _06497_ sky130_fd_sc_hd__nor3_1
XFILLER_0_77_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07143__A net1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13849_ _06418_ _06419_ VGND VGND VPWR VPWR _06421_ sky130_fd_sc_hd__xor2_1
XFILLER_0_9_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13799__B _02189_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07370_ _03400_ _03411_ VGND VGND VPWR VPWR _03422_ sky130_fd_sc_hd__and2b_1
XFILLER_0_85_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09040_ _01155_ _01156_ _01152_ _01154_ VGND VGND VPWR VPWR _01158_ sky130_fd_sc_hd__a211o_1
XFILLER_0_115_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09412__A1 _04510_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09412__B2 _00661_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap132 _06562_ VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__buf_1
Xmax_cap143 _01731_ VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09942_ _02109_ _02144_ VGND VGND VPWR VPWR _02145_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_111_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12224__A _00783_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10670__C _02849_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09873_ _02062_ _02067_ VGND VGND VPWR VPWR _02069_ sky130_fd_sc_hd__nand2_1
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08824_ _00919_ _00920_ VGND VGND VPWR VPWR _00921_ sky130_fd_sc_hd__and2b_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12878__B _01369_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08755_ _06637_ _00843_ _00845_ VGND VGND VPWR VPWR _00846_ sky130_fd_sc_hd__and3_1
XTAP_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07706_ _00880_ net64 VGND VGND VPWR VPWR _06835_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08686_ _05577_ _04048_ VGND VGND VPWR VPWR _00771_ sky130_fd_sc_hd__nand2_1
XTAP_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07637_ _05654_ _06329_ VGND VGND VPWR VPWR _06340_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07568_ _01405_ _05588_ VGND VGND VPWR VPWR _05599_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11589__A2 _01957_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09307_ _01319_ _01322_ VGND VGND VPWR VPWR _01450_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07499_ _04345_ _04356_ _04829_ VGND VGND VPWR VPWR _04840_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_91_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09238_ _01072_ _01078_ _01374_ VGND VGND VPWR VPWR _01375_ sky130_fd_sc_hd__and3_1
XFILLER_0_51_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09169_ _01187_ _01227_ _01297_ VGND VGND VPWR VPWR _01299_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_32_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11200_ _03525_ _03439_ VGND VGND VPWR VPWR _03526_ sky130_fd_sc_hd__nor2_2
XANTENNA__10013__A2 _00458_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12180_ _03582_ _03583_ VGND VGND VPWR VPWR _04603_ sky130_fd_sc_hd__or2_2
XANTENNA__11957__B _00138_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08612__A _06428_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07965__A1 _01120_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11131_ _03250_ _03449_ VGND VGND VPWR VPWR _03450_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11676__C _00755_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11062_ _03332_ _03321_ _03331_ VGND VGND VPWR VPWR _03374_ sky130_fd_sc_hd__nor3_1
X_10013_ _03015_ _00458_ _00608_ _00388_ VGND VGND VPWR VPWR _02223_ sky130_fd_sc_hd__a22o_1
XFILLER_0_25_16 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09162__B _02280_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11964_ _04292_ _04294_ _04364_ VGND VGND VPWR VPWR _04365_ sky130_fd_sc_hd__o21a_1
X_13703_ _06243_ _06247_ _06249_ VGND VGND VPWR VPWR _06260_ sky130_fd_sc_hd__nor3_1
X_10915_ _03209_ _03211_ VGND VGND VPWR VPWR _03212_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11895_ _04232_ _04251_ _04288_ VGND VGND VPWR VPWR _04289_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_129_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output109_A net109 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11029__A1 _00158_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13634_ _06181_ _06082_ _06183_ _06081_ VGND VGND VPWR VPWR _06184_ sky130_fd_sc_hd__a22o_1
X_10846_ _03124_ _03134_ _03135_ VGND VGND VPWR VPWR _03137_ sky130_fd_sc_hd__o21a_1
XFILLER_0_41_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13565_ _06106_ _06107_ VGND VGND VPWR VPWR _06108_ sky130_fd_sc_hd__or2_1
XFILLER_0_82_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10777_ _02116_ _02149_ _02723_ _02727_ VGND VGND VPWR VPWR _03061_ sky130_fd_sc_hd__and4_1
XFILLER_0_54_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12516_ _04970_ _04971_ VGND VGND VPWR VPWR _04973_ sky130_fd_sc_hd__and2b_1
XFILLER_0_81_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07653__B1 _06483_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13496_ _01415_ _03697_ _06020_ _06019_ VGND VGND VPWR VPWR _06033_ sky130_fd_sc_hd__a31o_1
XFILLER_0_14_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08225__C _00112_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12447_ _04886_ _04887_ VGND VGND VPWR VPWR _04897_ sky130_fd_sc_hd__xor2_1
XFILLER_0_140_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_output90_A net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10004__A2 _00612_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07405__B1 _03718_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08522__A _02007_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12378_ _04812_ _04820_ VGND VGND VPWR VPWR _04821_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10771__B _06461_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14117_ _06654_ _06713_ VGND VGND VPWR VPWR _06714_ sky130_fd_sc_hd__and2_1
X_11329_ _03640_ _03663_ VGND VGND VPWR VPWR _03668_ sky130_fd_sc_hd__xnor2_2
XANTENNA__07783__D _02960_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07138__A _00869_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14048_ _06639_ _06577_ _06630_ _06585_ VGND VGND VPWR VPWR _06640_ sky130_fd_sc_hd__a31o_1
X_08540_ _04268_ _04026_ _00446_ _00445_ VGND VGND VPWR VPWR _00611_ sky130_fd_sc_hd__a31oi_2
X_08471_ _00534_ _00535_ VGND VGND VPWR VPWR _00536_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_106_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08684__A2 _04015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07422_ _03839_ _03971_ VGND VGND VPWR VPWR _03993_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07353_ _01164_ _02609_ _02598_ VGND VGND VPWR VPWR _03235_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_17_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12219__A _00459_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08416__B _00003_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07284_ _02456_ _02467_ VGND VGND VPWR VPWR _02478_ sky130_fd_sc_hd__nand2_1
XFILLER_0_143_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09023_ _03543_ _00298_ _01138_ VGND VGND VPWR VPWR _01139_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_142_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11991__A2 _01958_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09247__B _02719_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07693__D _06821_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10951__B1 _01505_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09925_ _02124_ _02125_ VGND VGND VPWR VPWR _02126_ sky130_fd_sc_hd__or2b_1
X_09856_ _02045_ _02050_ VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__xnor2_1
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08807_ _00900_ _00902_ VGND VGND VPWR VPWR _00903_ sky130_fd_sc_hd__and2b_1
XFILLER_0_147_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09787_ _01818_ _01975_ VGND VGND VPWR VPWR _01976_ sky130_fd_sc_hd__xor2_1
XTAP_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08738_ _06885_ _00293_ VGND VGND VPWR VPWR _00828_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08669_ _05731_ net60 net8 net9 VGND VGND VPWR VPWR _00752_ sky130_fd_sc_hd__and4_1
XTAP_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10700_ _02963_ _02962_ VGND VGND VPWR VPWR _02976_ sky130_fd_sc_hd__and2b_1
XTAP_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12208__B1 _02135_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11680_ _04051_ _04052_ VGND VGND VPWR VPWR _04053_ sky130_fd_sc_hd__nor2_1
XTAP_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10232__A2_N _02459_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10856__B _02857_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10631_ _02810_ _02899_ VGND VGND VPWR VPWR _02900_ sky130_fd_sc_hd__xor2_1
XFILLER_0_107_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13350_ _05871_ _05872_ VGND VGND VPWR VPWR _05873_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10562_ _02821_ _02823_ VGND VGND VPWR VPWR _02824_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12301_ _04733_ _04735_ VGND VGND VPWR VPWR _04736_ sky130_fd_sc_hd__xor2_2
XFILLER_0_122_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13281_ _05598_ _05735_ _05803_ VGND VGND VPWR VPWR _05804_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_134_686 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10493_ _02247_ _02721_ VGND VGND VPWR VPWR _02748_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12232_ _04656_ _04658_ VGND VGND VPWR VPWR _04660_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12163_ _04583_ VGND VGND VPWR VPWR _04584_ sky130_fd_sc_hd__inv_2
XANTENNA__08060__B1 _06733_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08061__B _06744_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11114_ _02578_ _02545_ VGND VGND VPWR VPWR _03431_ sky130_fd_sc_hd__or2b_1
X_12094_ _04436_ _04439_ _04507_ VGND VGND VPWR VPWR _04508_ sky130_fd_sc_hd__o21a_1
X_11045_ _03353_ _03354_ VGND VGND VPWR VPWR _03355_ sky130_fd_sc_hd__and2_1
XFILLER_0_36_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09604__C _00414_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12996_ _05498_ _05499_ VGND VGND VPWR VPWR _05501_ sky130_fd_sc_hd__nand2_4
XFILLER_0_98_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11947_ _04274_ _04276_ VGND VGND VPWR VPWR _04347_ sky130_fd_sc_hd__and2_1
XANTENNA__07124__C net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11878_ _04269_ _04270_ VGND VGND VPWR VPWR _04271_ sky130_fd_sc_hd__and2_1
XFILLER_0_74_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13617_ _06163_ _06165_ VGND VGND VPWR VPWR _06166_ sky130_fd_sc_hd__and2b_1
X_10829_ _01350_ _02728_ _03117_ VGND VGND VPWR VPWR _03118_ sky130_fd_sc_hd__and3_1
XANTENNA__08418__A2 _00003_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11422__A1 _07004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13548_ _06084_ _06057_ _06088_ VGND VGND VPWR VPWR _06090_ sky130_fd_sc_hd__o21a_1
XFILLER_0_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_642 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12981__B _05483_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13479_ _06012_ VGND VGND VPWR VPWR _06014_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07929__A1 _00672_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12205__C _01953_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07971_ _00008_ _00013_ VGND VGND VPWR VPWR _00015_ sky130_fd_sc_hd__and2_1
XFILLER_0_10_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09710_ _01665_ _01669_ _01666_ VGND VGND VPWR VPWR _01891_ sky130_fd_sc_hd__o21ba_1
X_09641_ _01814_ _01815_ VGND VGND VPWR VPWR _01816_ sky130_fd_sc_hd__xnor2_1
X_09572_ _01739_ _01321_ VGND VGND VPWR VPWR _01740_ sky130_fd_sc_hd__and2b_1
XFILLER_0_93_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_846 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08523_ _00590_ _00591_ VGND VGND VPWR VPWR _00592_ sky130_fd_sc_hd__and2_1
XFILLER_0_77_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08454_ _00291_ _00302_ _00318_ VGND VGND VPWR VPWR _00517_ sky130_fd_sc_hd__o21a_1
XFILLER_0_77_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07331__A _02982_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07405_ _01394_ _03685_ _03718_ _01470_ VGND VGND VPWR VPWR _03806_ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08385_ _04279_ _04257_ VGND VGND VPWR VPWR _00441_ sky130_fd_sc_hd__or2b_1
XFILLER_0_147_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07336_ _03026_ _03037_ VGND VGND VPWR VPWR _03048_ sky130_fd_sc_hd__nor2_1
XANTENNA__11413__A1 _00268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11413__B2 _06733_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12891__B _02134_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07267_ _01799_ _01700_ _01788_ VGND VGND VPWR VPWR _02291_ sky130_fd_sc_hd__and3_1
XANTENNA__10692__A _00094_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11003__D _00959_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09006_ _01013_ _01016_ VGND VGND VPWR VPWR _01121_ sky130_fd_sc_hd__and2b_1
XFILLER_0_104_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07198_ _01492_ _01525_ VGND VGND VPWR VPWR _01536_ sky130_fd_sc_hd__or2b_4
XFILLER_0_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08593__A1 _06494_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09908_ _02106_ _02107_ VGND VGND VPWR VPWR _02108_ sky130_fd_sc_hd__xnor2_2
XANTENNA__07506__A _04906_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09839_ _01773_ _01806_ _02032_ VGND VGND VPWR VPWR _02033_ sky130_fd_sc_hd__a21o_1
XANTENNA__11028__A net6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12850_ _05266_ _05338_ _05339_ VGND VGND VPWR VPWR _05340_ sky130_fd_sc_hd__a21o_1
XFILLER_0_69_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11801_ _02674_ _02672_ VGND VGND VPWR VPWR _04186_ sky130_fd_sc_hd__or2b_1
XTAP_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12781_ _02305_ _05091_ _05263_ VGND VGND VPWR VPWR _05264_ sky130_fd_sc_hd__a21bo_1
XTAP_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11732_ _04076_ _02627_ _04077_ VGND VGND VPWR VPWR _04110_ sky130_fd_sc_hd__a21oi_1
XTAP_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08337__A _00389_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10586__B _04928_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07241__A _01996_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11663_ _00258_ _00414_ _00574_ _06765_ VGND VGND VPWR VPWR _04034_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13402_ _05397_ _05928_ VGND VGND VPWR VPWR _05930_ sky130_fd_sc_hd__or2_1
XFILLER_0_126_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10614_ _02878_ _02880_ VGND VGND VPWR VPWR _02881_ sky130_fd_sc_hd__or2b_1
XANTENNA__11404__A1 _00004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11594_ _03946_ _03957_ VGND VGND VPWR VPWR _03958_ sky130_fd_sc_hd__xor2_1
XFILLER_0_36_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13333_ _05325_ _05332_ VGND VGND VPWR VPWR _05854_ sky130_fd_sc_hd__nand2_1
X_10545_ _02801_ _02804_ VGND VGND VPWR VPWR _02805_ sky130_fd_sc_hd__or2b_1
XFILLER_0_52_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13264_ _05507_ _05524_ _05563_ VGND VGND VPWR VPWR _05788_ sky130_fd_sc_hd__and3_1
XANTENNA__08072__A _01350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10476_ _02728_ VGND VGND VPWR VPWR _02730_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__12306__B _01780_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12215_ _04639_ _03750_ _00458_ _04640_ VGND VGND VPWR VPWR _04641_ sky130_fd_sc_hd__and4b_1
X_13195_ _05717_ _05718_ VGND VGND VPWR VPWR _05719_ sky130_fd_sc_hd__nand2_1
X_12146_ _04557_ _04562_ _04564_ VGND VGND VPWR VPWR _04566_ sky130_fd_sc_hd__nor3_2
XFILLER_0_20_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12077_ _04487_ _04402_ _04489_ VGND VGND VPWR VPWR _04490_ sky130_fd_sc_hd__o21a_1
XFILLER_0_47_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11028_ net6 _04851_ _00780_ _00777_ VGND VGND VPWR VPWR _03337_ sky130_fd_sc_hd__and4_1
XANTENNA__10143__A1 _04862_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10143__B2 _04873_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11880__B _00670_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12979_ _04581_ _04584_ _04580_ _04486_ _05481_ VGND VGND VPWR VPWR _05482_ sky130_fd_sc_hd__a311oi_4
XANTENNA__10777__A _02116_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10496__B _00526_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08170_ _00211_ _00213_ VGND VGND VPWR VPWR _00214_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_103_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07121_ _00617_ _00683_ VGND VGND VPWR VPWR _00694_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13600__B _03783_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput101 net101 VGND VGND VPWR VPWR prod[42] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput112 net112 VGND VGND VPWR VPWR prod[52] sky130_fd_sc_hd__clkbuf_4
XANTENNA__08413__C _07010_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput123 net123 VGND VGND VPWR VPWR prod[62] sky130_fd_sc_hd__buf_4
XFILLER_0_11_632 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07954_ _06985_ _07000_ _07082_ VGND VGND VPWR VPWR _07083_ sky130_fd_sc_hd__o21a_1
XFILLER_0_49_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07326__A _00464_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07885_ _01120_ net37 VGND VGND VPWR VPWR _07014_ sky130_fd_sc_hd__nand2_1
X_09624_ _01573_ _01595_ VGND VGND VPWR VPWR _01797_ sky130_fd_sc_hd__or2_1
XANTENNA__09541__A _04598_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09555_ _01720_ _01485_ VGND VGND VPWR VPWR _01721_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08506_ _00572_ VGND VGND VPWR VPWR _00574_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_78_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09486_ _01644_ VGND VGND VPWR VPWR _01646_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07302__A2 _00672_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08437_ _05456_ _04895_ _00498_ VGND VGND VPWR VPWR _00499_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_108_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08368_ net9 VGND VGND VPWR VPWR _00423_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_135_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_510 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07319_ _00858_ _02850_ _02828_ _01853_ VGND VGND VPWR VPWR _02861_ sky130_fd_sc_hd__o211a_1
XFILLER_0_34_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08299_ _00251_ _00347_ VGND VGND VPWR VPWR _00348_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_6_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12407__A _00373_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10330_ _05027_ net40 _02369_ _02366_ VGND VGND VPWR VPWR _02570_ sky130_fd_sc_hd__a31o_1
XFILLER_0_33_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08015__B1 net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11030__B net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10261_ _01640_ _02046_ _02492_ _02494_ VGND VGND VPWR VPWR _02495_ sky130_fd_sc_hd__a31o_1
XFILLER_0_131_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12000_ _03990_ _03992_ VGND VGND VPWR VPWR _04405_ sky130_fd_sc_hd__and2_1
X_10192_ _02079_ _02417_ VGND VGND VPWR VPWR _02419_ sky130_fd_sc_hd__nand2_1
XANTENNA__14060__C _02743_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13311__A1 _05786_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13951_ _06521_ _06532_ VGND VGND VPWR VPWR _06533_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_17_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12902_ _05380_ _05396_ VGND VGND VPWR VPWR _05397_ sky130_fd_sc_hd__nand2_1
X_13882_ _06456_ VGND VGND VPWR VPWR _06457_ sky130_fd_sc_hd__inv_2
XANTENNA__12796__B _00392_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12833_ _05299_ _05301_ VGND VGND VPWR VPWR _05321_ sky130_fd_sc_hd__or2b_1
XTAP_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12764_ _05243_ _05244_ VGND VGND VPWR VPWR _05245_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11715_ _04089_ _04090_ VGND VGND VPWR VPWR _04091_ sky130_fd_sc_hd__nor2_1
XTAP_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12695_ _05161_ _05165_ _05168_ VGND VGND VPWR VPWR _05169_ sky130_fd_sc_hd__o21ba_1
XTAP_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_860 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11646_ _02249_ _04014_ VGND VGND VPWR VPWR _04016_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput14 a[21] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_4
Xinput25 a[31] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__buf_1
XANTENNA__13420__B _01181_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput36 b[12] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_4
X_11577_ _03909_ _03939_ VGND VGND VPWR VPWR _03940_ sky130_fd_sc_hd__xnor2_1
Xinput47 b[22] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__buf_4
XFILLER_0_40_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08514__B _01405_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput58 b[3] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__buf_8
XFILLER_0_52_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13316_ _05811_ _05835_ VGND VGND VPWR VPWR _05838_ sky130_fd_sc_hd__nor2_1
X_10528_ _02779_ _02786_ VGND VGND VPWR VPWR _02787_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13247_ _05757_ _05768_ _05769_ _02717_ _05772_ VGND VGND VPWR VPWR _05773_ sky130_fd_sc_hd__a221oi_4
XFILLER_0_0_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10459_ _02709_ _02710_ _02487_ VGND VGND VPWR VPWR _02712_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_440 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12353__A2 _00605_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13178_ _04403_ _04454_ VGND VGND VPWR VPWR _05701_ sky130_fd_sc_hd__nand2_1
X_12129_ _04541_ _04544_ VGND VGND VPWR VPWR _04547_ sky130_fd_sc_hd__nor2_1
X_07670_ _06340_ _06384_ _06604_ VGND VGND VPWR VPWR _06701_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_74_89 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09361__A _01383_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09340_ _01484_ _01485_ VGND VGND VPWR VPWR _01486_ sky130_fd_sc_hd__nand2_2
XANTENNA__10419__A2 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09271_ _01410_ VGND VGND VPWR VPWR _01411_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_90_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08222_ _00260_ _00265_ VGND VGND VPWR VPWR _00266_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_117_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08705__A _00431_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08153_ _06889_ _06888_ VGND VGND VPWR VPWR _00197_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07104_ _00497_ VGND VGND VPWR VPWR _00508_ sky130_fd_sc_hd__buf_4
XFILLER_0_43_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08084_ _00032_ _00127_ VGND VGND VPWR VPWR _00128_ sky130_fd_sc_hd__and2_1
XFILLER_0_70_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08440__A _02018_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13058__A _00381_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08986_ _01083_ _01097_ VGND VGND VPWR VPWR _01099_ sky130_fd_sc_hd__nand2_1
X_07937_ _07057_ _07064_ VGND VGND VPWR VPWR _07066_ sky130_fd_sc_hd__or2_1
XANTENNA__10107__A1 _05742_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10107__B2 _00628_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07868_ _06989_ _06995_ _06996_ VGND VGND VPWR VPWR _06997_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_3_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07523__A2 _00355_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08720__A1 _03532_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09271__A _01410_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08720__B2 _00121_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09607_ _01776_ _01778_ VGND VGND VPWR VPWR _01779_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07799_ _06926_ _06927_ VGND VGND VPWR VPWR _06928_ sky130_fd_sc_hd__nand2_2
XFILLER_0_97_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09538_ _01701_ _01702_ VGND VGND VPWR VPWR _01703_ sky130_fd_sc_hd__xor2_1
XANTENNA__07503__B _00311_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09276__A2 _01062_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09469_ _01626_ _01560_ _01561_ VGND VGND VPWR VPWR _01628_ sky130_fd_sc_hd__nor3_1
XFILLER_0_54_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11500_ _03721_ _03854_ VGND VGND VPWR VPWR _03855_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10830__A2 net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12480_ _04817_ _04819_ VGND VGND VPWR VPWR _04933_ sky130_fd_sc_hd__and2_1
XFILLER_0_108_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11431_ _03769_ _03771_ VGND VGND VPWR VPWR _03779_ sky130_fd_sc_hd__nand2_1
XFILLER_0_80_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14150_ _06747_ _06748_ VGND VGND VPWR VPWR _06749_ sky130_fd_sc_hd__nand2_1
XANTENNA__09984__B1 _02190_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11362_ _02246_ _03687_ _03684_ _02249_ VGND VGND VPWR VPWR _03703_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13101_ _04551_ _04531_ VGND VGND VPWR VPWR _05616_ sky130_fd_sc_hd__and2_1
XFILLER_0_21_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10313_ _05203_ _00604_ VGND VGND VPWR VPWR _02551_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14081_ _06673_ _06674_ VGND VGND VPWR VPWR _06675_ sky130_fd_sc_hd__nand2_1
X_11293_ _02757_ _02788_ VGND VGND VPWR VPWR _03628_ sky130_fd_sc_hd__and2_1
X_13032_ _05532_ _05539_ VGND VGND VPWR VPWR _05540_ sky130_fd_sc_hd__or2_1
X_10244_ _02473_ _02475_ VGND VGND VPWR VPWR _02476_ sky130_fd_sc_hd__nor2_1
XANTENNA__11695__B _06875_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09446__A _02335_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08350__A _00464_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09200__A2 _00144_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10175_ _00101_ _03685_ _03718_ net37 VGND VGND VPWR VPWR _02400_ sky130_fd_sc_hd__a22o_1
XANTENNA__12022__D _03679_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13934_ _06511_ _06513_ VGND VGND VPWR VPWR _06514_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07514__A2 _04851_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09181__A _00654_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13048__B1 _00393_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13865_ _06422_ _06437_ VGND VGND VPWR VPWR _06438_ sky130_fd_sc_hd__and2_1
XANTENNA__08509__B _00311_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13599__A1 _01061_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12816_ _05299_ _05301_ VGND VGND VPWR VPWR _05303_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13599__B2 _02856_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13796_ _06311_ _06359_ _06361_ VGND VGND VPWR VPWR _06363_ sky130_fd_sc_hd__o21a_1
XFILLER_0_146_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12747_ _00379_ _03678_ VGND VGND VPWR VPWR _05227_ sky130_fd_sc_hd__nand2_1
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10821__A2 net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12678_ _05133_ _05134_ VGND VGND VPWR VPWR _05151_ sky130_fd_sc_hd__xor2_1
XANTENNA__10774__B _02168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11629_ _03983_ _03994_ _03996_ VGND VGND VPWR VPWR _03997_ sky130_fd_sc_hd__a21oi_2
XANTENNA__12023__A1 _06626_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12023__B2 _06450_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09356__A _01369_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08840_ _00740_ _00937_ _00938_ VGND VGND VPWR VPWR _00939_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_85_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12213__C _01179_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08771_ _00696_ _00699_ _00863_ VGND VGND VPWR VPWR _00864_ sky130_fd_sc_hd__nor3_1
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10014__B _02971_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13826__A2 _03683_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07722_ _06790_ _06850_ VGND VGND VPWR VPWR _06851_ sky130_fd_sc_hd__nor2_1
X_07653_ _06428_ _06472_ _06483_ _06439_ VGND VGND VPWR VPWR _06516_ sky130_fd_sc_hd__a22o_1
X_07584_ _05753_ _05761_ _00901_ _02664_ VGND VGND VPWR VPWR _05771_ sky130_fd_sc_hd__and4b_1
XFILLER_0_47_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09323_ _01465_ _01466_ VGND VGND VPWR VPWR _01467_ sky130_fd_sc_hd__and2_1
XFILLER_0_87_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09254_ _01381_ _01095_ _01390_ VGND VGND VPWR VPWR _01392_ sky130_fd_sc_hd__nor3_1
XANTENNA__12875__A1_N _01180_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08205_ _00206_ _00242_ _00245_ _00246_ _00248_ VGND VGND VPWR VPWR _00249_ sky130_fd_sc_hd__o32ai_4
XFILLER_0_106_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09185_ _01313_ _01315_ VGND VGND VPWR VPWR _01316_ sky130_fd_sc_hd__and2_1
XFILLER_0_50_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08136_ _00178_ _00083_ _00179_ VGND VGND VPWR VPWR _00180_ sky130_fd_sc_hd__nor3_2
XFILLER_0_71_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_524 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08067_ _00009_ _00010_ _00011_ VGND VGND VPWR VPWR _00111_ sky130_fd_sc_hd__and3_1
XFILLER_0_113_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12317__A2 _02088_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12404__B _01272_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08969_ _01071_ _01079_ VGND VGND VPWR VPWR _01080_ sky130_fd_sc_hd__xor2_1
X_11980_ _04316_ _04212_ _04317_ VGND VGND VPWR VPWR _04383_ sky130_fd_sc_hd__or3_2
XANTENNA__10859__B _01410_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10931_ _02520_ _03226_ _03228_ VGND VGND VPWR VPWR _03230_ sky130_fd_sc_hd__o21a_1
XFILLER_0_98_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13650_ _06195_ _06200_ _06191_ VGND VGND VPWR VPWR _06202_ sky130_fd_sc_hd__a21oi_1
X_10862_ _03149_ _03152_ _03153_ VGND VGND VPWR VPWR _03154_ sky130_fd_sc_hd__and3_1
XFILLER_0_14_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12601_ _05050_ _05048_ VGND VGND VPWR VPWR _05066_ sky130_fd_sc_hd__and2b_1
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13581_ _06122_ _06125_ VGND VGND VPWR VPWR _06126_ sky130_fd_sc_hd__or2_1
XFILLER_0_137_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10793_ _06937_ _02758_ _03075_ _03076_ VGND VGND VPWR VPWR _03078_ sky130_fd_sc_hd__a22oi_1
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13251__A _05776_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12532_ _04930_ _04988_ _04989_ VGND VGND VPWR VPWR _04990_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_94_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08345__A _00352_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10594__B _00310_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08209__B1 _00100_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07680__A1 net1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12463_ _04812_ _04820_ VGND VGND VPWR VPWR _04914_ sky130_fd_sc_hd__or2_1
XANTENNA__12005__A1 _00843_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07680__B2 net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12005__B2 _00844_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14202_ _02938_ _02927_ VGND VGND VPWR VPWR _06794_ sky130_fd_sc_hd__and2b_2
XFILLER_0_50_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11414_ _03758_ _03759_ VGND VGND VPWR VPWR _03760_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12394_ _00778_ _00413_ _00571_ _00782_ VGND VGND VPWR VPWR _04838_ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_395 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14133_ _06077_ _04013_ _06705_ _06704_ VGND VGND VPWR VPWR _06730_ sky130_fd_sc_hd__a31o_1
X_11345_ _03683_ VGND VGND VPWR VPWR _03684_ sky130_fd_sc_hd__buf_2
XFILLER_0_1_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14064_ _06654_ _06655_ VGND VGND VPWR VPWR _06656_ sky130_fd_sc_hd__or2_1
X_11276_ _03604_ _03607_ VGND VGND VPWR VPWR _03610_ sky130_fd_sc_hd__or2_1
XANTENNA__12314__B _01780_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13015_ _05520_ _05495_ VGND VGND VPWR VPWR _05521_ sky130_fd_sc_hd__xnor2_2
X_10227_ _02447_ _02457_ VGND VGND VPWR VPWR _02458_ sky130_fd_sc_hd__xor2_1
XFILLER_0_146_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10158_ _02378_ _02381_ VGND VGND VPWR VPWR _02382_ sky130_fd_sc_hd__or2_2
XFILLER_0_55_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10089_ _02158_ VGND VGND VPWR VPWR _02306_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__07424__A net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13917_ _06363_ _06495_ VGND VGND VPWR VPWR _06496_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13848_ _06418_ _06419_ VGND VGND VPWR VPWR _06420_ sky130_fd_sc_hd__nand2_1
XFILLER_0_147_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13441__B1 _02735_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13779_ _06332_ _06333_ VGND VGND VPWR VPWR _06344_ sky130_fd_sc_hd__nor2_1
XANTENNA__13799__C _03686_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08255__A _00157_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09412__A2 _01177_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_cap133 net134 VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap144 _04299_ VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__buf_1
XANTENNA__12505__A _04037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09941_ _02142_ _02143_ VGND VGND VPWR VPWR _02144_ sky130_fd_sc_hd__or2_1
XFILLER_0_40_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12224__B _00778_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10670__D _02304_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_798 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09872_ _02062_ _02067_ VGND VGND VPWR VPWR _02068_ sky130_fd_sc_hd__nor2_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08823_ _01044_ net8 _03718_ _05731_ VGND VGND VPWR VPWR _00920_ sky130_fd_sc_hd__a22o_1
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13336__A _00914_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12878__C _01248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08754_ _06937_ _00844_ VGND VGND VPWR VPWR _00845_ sky130_fd_sc_hd__nand2_1
XTAP_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07705_ _06802_ _06797_ VGND VGND VPWR VPWR _06834_ sky130_fd_sc_hd__or2b_1
XTAP_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08685_ _00767_ _00768_ VGND VGND VPWR VPWR _00769_ sky130_fd_sc_hd__and2b_1
XFILLER_0_95_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07636_ _05934_ _06318_ VGND VGND VPWR VPWR _06329_ sky130_fd_sc_hd__xnor2_1
XTAP_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07567_ _05577_ VGND VGND VPWR VPWR _05588_ sky130_fd_sc_hd__buf_4
XFILLER_0_48_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09306_ _01318_ _01323_ VGND VGND VPWR VPWR _01449_ sky130_fd_sc_hd__and2b_1
XFILLER_0_119_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07498_ _04587_ _04818_ VGND VGND VPWR VPWR _04829_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_118_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09237_ _01367_ _01373_ VGND VGND VPWR VPWR _01374_ sky130_fd_sc_hd__xor2_1
XFILLER_0_17_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09168_ _01187_ _01227_ _01297_ VGND VGND VPWR VPWR _01298_ sky130_fd_sc_hd__and3_1
XFILLER_0_133_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08119_ _00066_ _00067_ _00064_ VGND VGND VPWR VPWR _00163_ sky130_fd_sc_hd__o21ba_1
XANTENNA__08611__B1 _00310_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09099_ _01221_ _01222_ VGND VGND VPWR VPWR _01223_ sky130_fd_sc_hd__nor2_1
XANTENNA__11957__C _02134_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08612__B _06439_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07965__A2 net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11130_ _03305_ _03447_ _03448_ VGND VGND VPWR VPWR _03449_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_101_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11676__D _01260_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11061_ _03289_ _03372_ VGND VGND VPWR VPWR _03373_ sky130_fd_sc_hd__nor2_1
XANTENNA__07178__B1 _01306_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10012_ _02220_ _02221_ VGND VGND VPWR VPWR _02222_ sky130_fd_sc_hd__xor2_2
XFILLER_0_99_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08193__B1_N _00208_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_332 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07244__A _02029_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_28 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11963_ _04362_ _04363_ VGND VGND VPWR VPWR _04364_ sky130_fd_sc_hd__nor2_1
XANTENNA__09162__C _00416_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10485__B1 _02737_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13702_ _06247_ _06257_ _06258_ VGND VGND VPWR VPWR _06259_ sky130_fd_sc_hd__or3_1
X_10914_ _03161_ _03210_ VGND VGND VPWR VPWR _03211_ sky130_fd_sc_hd__nor2_1
X_11894_ _04216_ _04231_ VGND VGND VPWR VPWR _04288_ sky130_fd_sc_hd__and2b_1
X_13633_ _06181_ _06182_ VGND VGND VPWR VPWR _06183_ sky130_fd_sc_hd__nand2_1
X_10845_ _03116_ _03118_ VGND VGND VPWR VPWR _03135_ sky130_fd_sc_hd__xor2_1
XANTENNA__11029__A2 _04037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13564_ _06074_ _04014_ _06104_ _06105_ VGND VGND VPWR VPWR _06107_ sky130_fd_sc_hd__and4_1
X_10776_ _02160_ _02723_ _02727_ _02116_ VGND VGND VPWR VPWR _03060_ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07653__A1 _06428_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12515_ _00374_ _04059_ _03707_ _03740_ VGND VGND VPWR VPWR _04971_ sky130_fd_sc_hd__and4_2
XFILLER_0_109_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13495_ _06017_ _06030_ VGND VGND VPWR VPWR _06031_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07653__B2 _06439_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07410__C net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08225__D _00268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12446_ _04893_ _04894_ VGND VGND VPWR VPWR _04896_ sky130_fd_sc_hd__nor2_1
XFILLER_0_140_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07405__B2 _01470_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12377_ _04817_ _04819_ VGND VGND VPWR VPWR _04820_ sky130_fd_sc_hd__nor2_1
XFILLER_0_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08522__B _02040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10771__C _02724_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output83_A net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14116_ _06673_ _06711_ VGND VGND VPWR VPWR _06713_ sky130_fd_sc_hd__xnor2_1
X_11328_ _03627_ _03666_ VGND VGND VPWR VPWR _03667_ sky130_fd_sc_hd__xnor2_2
X_14047_ net132 VGND VGND VPWR VPWR _06639_ sky130_fd_sc_hd__inv_2
X_11259_ _03570_ _03571_ VGND VGND VPWR VPWR _03591_ sky130_fd_sc_hd__nand2_1
XANTENNA__09634__A _01197_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08470_ _03532_ _00151_ VGND VGND VPWR VPWR _00535_ sky130_fd_sc_hd__nand2_1
XFILLER_0_106_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07421_ _03839_ _03971_ VGND VGND VPWR VPWR _03982_ sky130_fd_sc_hd__nor2_1
XFILLER_0_106_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07892__A1 _00541_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07352_ _03202_ _03213_ VGND VGND VPWR VPWR _03224_ sky130_fd_sc_hd__or2_4
XFILLER_0_116_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12219__B _00608_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07283_ _02259_ VGND VGND VPWR VPWR _02467_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_45_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09022_ _01135_ _01136_ _01137_ VGND VGND VPWR VPWR _01138_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_115_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12235__A _00783_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07329__A _02960_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10951__A1 _00143_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10951__B2 _04906_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09924_ _02114_ _02123_ VGND VGND VPWR VPWR _02125_ sky130_fd_sc_hd__nand2_1
XFILLER_0_111_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09855_ _01640_ _02046_ _02049_ VGND VGND VPWR VPWR _02050_ sky130_fd_sc_hd__a21oi_1
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08806_ _03850_ net13 _00730_ _01394_ VGND VGND VPWR VPWR _00902_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09786_ _01972_ _01973_ VGND VGND VPWR VPWR _01975_ sky130_fd_sc_hd__and2b_1
XTAP_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08737_ _00258_ _00656_ _00826_ VGND VGND VPWR VPWR _00827_ sky130_fd_sc_hd__a21bo_1
XTAP_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08668_ _00747_ _00750_ VGND VGND VPWR VPWR _00751_ sky130_fd_sc_hd__xnor2_2
XTAP_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12208__A1 _01518_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07619_ _06131_ _02883_ _02445_ _03477_ VGND VGND VPWR VPWR _06142_ sky130_fd_sc_hd__nand4b_4
XTAP_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08599_ _00479_ _00675_ VGND VGND VPWR VPWR _00676_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10630_ _00818_ _02731_ _02898_ VGND VGND VPWR VPWR _02899_ sky130_fd_sc_hd__and3_1
XFILLER_0_76_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10561_ _02818_ _02822_ VGND VGND VPWR VPWR _02823_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_91_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12300_ _02190_ _02426_ _04734_ VGND VGND VPWR VPWR _04735_ sky130_fd_sc_hd__and3_1
XFILLER_0_133_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13280_ _05728_ _05730_ VGND VGND VPWR VPWR _05803_ sky130_fd_sc_hd__and2_1
XFILLER_0_63_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10492_ _02733_ _02732_ VGND VGND VPWR VPWR _02747_ sky130_fd_sc_hd__or2b_1
XFILLER_0_106_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12231_ _04656_ _04658_ VGND VGND VPWR VPWR _04659_ sky130_fd_sc_hd__nand2_1
XFILLER_0_133_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12162_ _04484_ _04582_ VGND VGND VPWR VPWR _04583_ sky130_fd_sc_hd__or2b_1
XANTENNA__08060__A1 _02105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08060__B2 _00650_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11113_ _03421_ _03429_ VGND VGND VPWR VPWR _03430_ sky130_fd_sc_hd__xnor2_1
X_12093_ _04505_ _04506_ VGND VGND VPWR VPWR _04507_ sky130_fd_sc_hd__nor2_1
X_11044_ _03346_ _03349_ VGND VGND VPWR VPWR _03354_ sky130_fd_sc_hd__xor2_1
XFILLER_0_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09604__D _00574_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output121_A net121 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12995_ _00381_ _02008_ _05497_ _05022_ VGND VGND VPWR VPWR _05499_ sky130_fd_sc_hd__a211o_1
XFILLER_0_86_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11946_ _04274_ _04276_ _04344_ VGND VGND VPWR VPWR _04346_ sky130_fd_sc_hd__and3_1
XFILLER_0_143_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07702__A net1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11877_ _04256_ _04267_ VGND VGND VPWR VPWR _04270_ sky130_fd_sc_hd__or2_1
X_13616_ _06140_ _06143_ VGND VGND VPWR VPWR _06165_ sky130_fd_sc_hd__xor2_1
X_10828_ _01383_ _02724_ VGND VGND VPWR VPWR _03117_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07626__A1 _05445_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13547_ _06084_ _06057_ _06088_ VGND VGND VPWR VPWR _06089_ sky130_fd_sc_hd__nor3_1
XANTENNA__08823__B1 _03718_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11422__A2 _03748_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10759_ _03038_ _03040_ VGND VGND VPWR VPWR _03041_ sky130_fd_sc_hd__nor2_1
XFILLER_0_70_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13478_ _06011_ _06012_ _01062_ _03684_ VGND VGND VPWR VPWR _06013_ sky130_fd_sc_hd__and4b_1
XFILLER_0_140_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12429_ _04761_ _04769_ VGND VGND VPWR VPWR _04877_ sky130_fd_sc_hd__xor2_1
XFILLER_0_124_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07929__A2 _05027_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07149__A net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07970_ _00008_ _00013_ VGND VGND VPWR VPWR _00014_ sky130_fd_sc_hd__nor2_1
XANTENNA__12205__D _02134_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09640_ _00311_ net20 VGND VGND VPWR VPWR _01815_ sky130_fd_sc_hd__nand2_1
X_09571_ _01450_ _01452_ _01455_ VGND VGND VPWR VPWR _01739_ sky130_fd_sc_hd__a21o_1
XFILLER_0_117_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08522_ _02007_ _02040_ _03707_ _00392_ VGND VGND VPWR VPWR _00591_ sky130_fd_sc_hd__nand4_4
XFILLER_0_78_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08708__A _04081_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08453_ _00513_ _00515_ VGND VGND VPWR VPWR _00516_ sky130_fd_sc_hd__or2_1
XFILLER_0_147_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07404_ _01394_ _01470_ _03685_ _03718_ VGND VGND VPWR VPWR _03795_ sky130_fd_sc_hd__and4_1
X_08384_ _02467_ _00381_ VGND VGND VPWR VPWR _00440_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07335_ _01470_ net33 _00355_ _02971_ VGND VGND VPWR VPWR _03037_ sky130_fd_sc_hd__and4_1
XFILLER_0_116_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11413__A2 _01178_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09539__A _00355_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07266_ _02040_ VGND VGND VPWR VPWR _02280_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_60_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10692__B _01411_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_143_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09005_ _06885_ _00294_ _01014_ VGND VGND VPWR VPWR _01119_ sky130_fd_sc_hd__and3_1
XFILLER_0_116_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07197_ _01284_ _00672_ _01503_ _01514_ VGND VGND VPWR VPWR _01525_ sky130_fd_sc_hd__a31o_1
XFILLER_0_103_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08593__A2 _00004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14180__A _02743_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09274__A _01413_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09907_ _02003_ _02005_ _02001_ VGND VGND VPWR VPWR _02107_ sky130_fd_sc_hd__a21o_1
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09838_ _01773_ _01806_ _01820_ VGND VGND VPWR VPWR _02032_ sky130_fd_sc_hd__o21a_1
XANTENNA__11028__B _04851_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09769_ _01955_ VGND VGND VPWR VPWR _01956_ sky130_fd_sc_hd__clkbuf_4
XTAP_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11800_ _04178_ _04184_ VGND VGND VPWR VPWR _04185_ sky130_fd_sc_hd__xor2_1
XTAP_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12780_ _00572_ _02849_ _02305_ _00414_ VGND VGND VPWR VPWR _05263_ sky130_fd_sc_hd__a22o_1
XTAP_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11731_ _02612_ _04108_ VGND VGND VPWR VPWR _04109_ sky130_fd_sc_hd__xnor2_1
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10586__C _02849_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11662_ _00258_ _06765_ _00414_ VGND VGND VPWR VPWR _04033_ sky130_fd_sc_hd__and3_1
X_13401_ _05397_ _05928_ VGND VGND VPWR VPWR _05929_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_850 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10613_ _02853_ _02879_ VGND VGND VPWR VPWR _02880_ sky130_fd_sc_hd__nand2_1
X_11593_ _03943_ _03944_ VGND VGND VPWR VPWR _03957_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11404__A2 _03748_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10544_ _00819_ _02169_ _02802_ _02803_ VGND VGND VPWR VPWR _02804_ sky130_fd_sc_hd__a31o_1
XFILLER_0_106_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13332_ _05362_ _05408_ VGND VGND VPWR VPWR _05853_ sky130_fd_sc_hd__and2b_1
XFILLER_0_91_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13263_ _05474_ _05490_ VGND VGND VPWR VPWR _05787_ sky130_fd_sc_hd__xnor2_4
X_10475_ _02727_ VGND VGND VPWR VPWR _02728_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08072__B _00113_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12214_ _01507_ _01179_ _01254_ _00605_ VGND VGND VPWR VPWR _04640_ sky130_fd_sc_hd__a22o_1
X_13194_ _05700_ _05704_ VGND VGND VPWR VPWR _05718_ sky130_fd_sc_hd__xor2_2
X_12145_ _04558_ _04561_ _04559_ _04563_ VGND VGND VPWR VPWR _04564_ sky130_fd_sc_hd__o31a_1
XFILLER_0_47_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12076_ _04452_ _04453_ VGND VGND VPWR VPWR _04489_ sky130_fd_sc_hd__nand2_1
XANTENNA__11219__A _00410_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11027_ _05027_ _00780_ _00777_ _04851_ VGND VGND VPWR VPWR _03336_ sky130_fd_sc_hd__a22o_1
XANTENNA__10143__A2 _00373_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11880__C _00915_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12978_ _04581_ _04584_ _04575_ VGND VGND VPWR VPWR _05481_ sky130_fd_sc_hd__and3_1
XANTENNA__10777__B _02149_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07432__A net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11929_ _04253_ _04322_ VGND VGND VPWR VPWR _04327_ sky130_fd_sc_hd__nor2_1
XANTENNA__10496__C _02735_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07120_ _00628_ _00650_ _00672_ _00300_ VGND VGND VPWR VPWR _00683_ sky130_fd_sc_hd__and4_1
XFILLER_0_55_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput102 net102 VGND VGND VPWR VPWR prod[43] sky130_fd_sc_hd__clkbuf_4
Xoutput113 net129 VGND VGND VPWR VPWR prod[53] sky130_fd_sc_hd__clkbuf_4
Xoutput124 net124 VGND VGND VPWR VPWR prod[63] sky130_fd_sc_hd__clkbuf_4
XANTENNA__08413__D _00101_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_644 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12513__A _04059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07953_ _07001_ _07081_ VGND VGND VPWR VPWR _07082_ sky130_fd_sc_hd__xnor2_2
X_07884_ _07011_ _07012_ VGND VGND VPWR VPWR _07013_ sky130_fd_sc_hd__nor2_1
XANTENNA__07326__B _00530_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09822__A _06821_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09623_ _01790_ _01795_ VGND VGND VPWR VPWR _01796_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10968__A _04862_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09541__B net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09554_ _01479_ _01719_ VGND VGND VPWR VPWR _01720_ sky130_fd_sc_hd__nand2_1
XANTENNA__11792__A1_N _02127_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08438__A _05456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08505_ _00571_ VGND VGND VPWR VPWR _00572_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_38_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09485_ _01631_ _01632_ VGND VGND VPWR VPWR _01644_ sky130_fd_sc_hd__or2_1
XANTENNA__09260__C _00605_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08436_ _05478_ _00142_ VGND VGND VPWR VPWR _00498_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08367_ _03850_ _04510_ net9 net10 VGND VGND VPWR VPWR _00422_ sky130_fd_sc_hd__and4_1
XFILLER_0_80_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07318_ _01219_ _01438_ _01842_ _01186_ VGND VGND VPWR VPWR _02850_ sky130_fd_sc_hd__o31a_1
XFILLER_0_34_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08263__A1 _02040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08298_ _00345_ _00346_ VGND VGND VPWR VPWR _00347_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08263__B2 _04917_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12407__B _00782_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07249_ _02072_ net184 VGND VGND VPWR VPWR _02094_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10260_ _02045_ _02049_ _02274_ _02493_ _02273_ VGND VGND VPWR VPWR _02494_ sky130_fd_sc_hd__a32o_1
XANTENNA__08015__A1 _01197_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08015__B2 _01208_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11030__C _00612_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10191_ _02079_ _02417_ VGND VGND VPWR VPWR _02418_ sky130_fd_sc_hd__or2_1
XANTENNA__07517__A _00300_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14060__D _02742_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13950_ _06523_ _06530_ _06531_ VGND VGND VPWR VPWR _06532_ sky130_fd_sc_hd__o21ba_2
X_12901_ _05394_ _05395_ VGND VGND VPWR VPWR _05396_ sky130_fd_sc_hd__and2_1
XFILLER_0_88_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13881_ _06454_ _06455_ VGND VGND VPWR VPWR _06456_ sky130_fd_sc_hd__and2_1
XANTENNA__12796__C _02168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12832_ _05295_ _05298_ VGND VGND VPWR VPWR _05320_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_110 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07252__A _00672_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12763_ _04647_ _05242_ VGND VGND VPWR VPWR _05244_ sky130_fd_sc_hd__and2b_1
XTAP_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11714_ _04088_ _04084_ _04085_ VGND VGND VPWR VPWR _04090_ sky130_fd_sc_hd__nor3_1
XTAP_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12694_ _05161_ _05165_ _05167_ VGND VGND VPWR VPWR _05168_ sky130_fd_sc_hd__a21boi_1
XTAP_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11645_ _03697_ VGND VGND VPWR VPWR _04014_ sky130_fd_sc_hd__buf_2
XFILLER_0_25_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput15 a[22] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__buf_4
XANTENNA__13420__C _01414_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput26 a[3] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_4
X_11576_ _00262_ _03748_ _03937_ VGND VGND VPWR VPWR _03939_ sky130_fd_sc_hd__and3_1
Xinput37 b[13] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_4
Xinput48 b[23] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08514__C _03773_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13315_ _05835_ VGND VGND VPWR VPWR _05836_ sky130_fd_sc_hd__inv_2
Xinput59 b[4] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__buf_4
XFILLER_0_134_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10527_ _02777_ _02778_ VGND VGND VPWR VPWR _02786_ sky130_fd_sc_hd__or2_1
XFILLER_0_107_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10118__A _06637_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13246_ _05592_ _05767_ _05770_ VGND VGND VPWR VPWR _05772_ sky130_fd_sc_hd__a21oi_2
X_10458_ _02487_ _02709_ _02710_ VGND VGND VPWR VPWR _02711_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08811__A _00300_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13177_ _03622_ _05699_ VGND VGND VPWR VPWR _05700_ sky130_fd_sc_hd__xnor2_2
X_10389_ _02399_ _02409_ VGND VGND VPWR VPWR _02635_ sky130_fd_sc_hd__nand2_1
XANTENNA__07427__A net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12128_ _04540_ _03955_ _04545_ VGND VGND VPWR VPWR _04546_ sky130_fd_sc_hd__mux2_2
XANTENNA__13148__B _05651_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12059_ _04469_ VGND VGND VPWR VPWR _04470_ sky130_fd_sc_hd__inv_2
XANTENNA__09361__B _01508_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09270_ net50 VGND VGND VPWR VPWR _01410_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_716 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08221_ _00120_ _00123_ _00261_ _00264_ VGND VGND VPWR VPWR _00265_ sky130_fd_sc_hd__a211o_2
XFILLER_0_118_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08705__B _04169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08152_ _06990_ _00195_ VGND VGND VPWR VPWR _00196_ sky130_fd_sc_hd__nor2_1
XANTENNA__11412__A _00114_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09442__B1 _00574_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07103_ _00486_ VGND VGND VPWR VPWR _00497_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_126_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11131__B _03449_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08083_ _00119_ _00126_ VGND VGND VPWR VPWR _00127_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_141_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_791 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09817__A _00530_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08440__B _00158_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07337__A _02018_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13058__B _00391_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08985_ _01095_ _01096_ VGND VGND VPWR VPWR _01097_ sky130_fd_sc_hd__nor2_1
XFILLER_0_139_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07936_ _07057_ _07064_ VGND VGND VPWR VPWR _07065_ sky130_fd_sc_hd__and2_1
XANTENNA__10107__A2 net50 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07867_ _06994_ _06991_ _06992_ VGND VGND VPWR VPWR _06996_ sky130_fd_sc_hd__and3_1
XFILLER_0_98_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08720__A2 _04895_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09606_ _03059_ _01600_ VGND VGND VPWR VPWR _01778_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07798_ _06924_ _06925_ _06923_ VGND VGND VPWR VPWR _06927_ sky130_fd_sc_hd__o21ai_1
X_09537_ _05192_ _04026_ VGND VGND VPWR VPWR _01702_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07503__C _04862_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09468_ _01560_ _01561_ _01626_ VGND VGND VPWR VPWR _01627_ sky130_fd_sc_hd__o21a_1
X_08419_ _00477_ _00478_ VGND VGND VPWR VPWR _00479_ sky130_fd_sc_hd__and2b_1
XFILLER_0_81_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09399_ _01549_ _01550_ VGND VGND VPWR VPWR _01551_ sky130_fd_sc_hd__xor2_1
XFILLER_0_46_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11430_ _03776_ _03777_ VGND VGND VPWR VPWR _03778_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11361_ _00843_ _00844_ _03687_ _03684_ VGND VGND VPWR VPWR _03702_ sky130_fd_sc_hd__and4_1
XANTENNA__09984__A1 _06637_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09984__B2 _06937_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_739 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13100_ _05612_ _05614_ VGND VGND VPWR VPWR _05615_ sky130_fd_sc_hd__and2_1
XFILLER_0_131_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10312_ _01369_ _02548_ _02549_ VGND VGND VPWR VPWR _02550_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_61_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14080_ _06661_ _06672_ VGND VGND VPWR VPWR _06674_ sky130_fd_sc_hd__or2_1
X_11292_ _02746_ _02790_ VGND VGND VPWR VPWR _03627_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_104_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13031_ _05536_ _05538_ VGND VGND VPWR VPWR _05539_ sky130_fd_sc_hd__or2_2
X_10243_ _02086_ _02108_ _02474_ VGND VGND VPWR VPWR _02475_ sky130_fd_sc_hd__o21ai_2
XANTENNA__09446__B _01601_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11695__C _01272_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08350__B _00381_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10174_ _02397_ _02398_ VGND VGND VPWR VPWR _02399_ sky130_fd_sc_hd__xnor2_2
X_13933_ _06482_ _06512_ VGND VGND VPWR VPWR _06513_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13048__A1 _00376_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10401__A _05445_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13864_ _05907_ _05911_ _06421_ VGND VGND VPWR VPWR _06437_ sky130_fd_sc_hd__or3_1
XANTENNA__08078__A _06461_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13048__B2 _00381_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08509__C _00413_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12815_ _05118_ _05129_ _05300_ VGND VGND VPWR VPWR _05301_ sky130_fd_sc_hd__a21o_1
XANTENNA__13599__A2 _03785_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13795_ _06290_ _06360_ VGND VGND VPWR VPWR _06361_ sky130_fd_sc_hd__nor2_1
XFILLER_0_57_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12746_ _00378_ _03681_ _04632_ _04630_ VGND VGND VPWR VPWR _05226_ sky130_fd_sc_hd__a31o_1
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12328__A _01066_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12677_ _05147_ _05149_ VGND VGND VPWR VPWR _05150_ sky130_fd_sc_hd__nand2_2
X_11628_ _03969_ _03995_ VGND VGND VPWR VPWR _03996_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12023__A2 _03683_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11559_ _00486_ _01960_ VGND VGND VPWR VPWR _03920_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09637__A _01744_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13229_ _05579_ _05755_ VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__xnor2_4
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07157__A _01076_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09075__C _01996_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12213__D _01254_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08770_ _00861_ _00862_ VGND VGND VPWR VPWR _00863_ sky130_fd_sc_hd__nor2_1
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10014__C net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07721_ _06829_ _06849_ VGND VGND VPWR VPWR _06850_ sky130_fd_sc_hd__xor2_2
XFILLER_0_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07652_ _06428_ _06450_ _06472_ _06494_ VGND VGND VPWR VPWR _06505_ sky130_fd_sc_hd__nand4_2
X_07583_ _05731_ _00628_ _05742_ _01000_ VGND VGND VPWR VPWR _05761_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09322_ _01447_ _01464_ VGND VGND VPWR VPWR _01466_ sky130_fd_sc_hd__or2_1
XANTENNA__08466__A1 _03543_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09253_ _01381_ _01095_ _01390_ VGND VGND VPWR VPWR _01391_ sky130_fd_sc_hd__o21a_1
XFILLER_0_35_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08204_ _00247_ VGND VGND VPWR VPWR _00248_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09184_ _01314_ VGND VGND VPWR VPWR _01315_ sky130_fd_sc_hd__inv_2
X_08135_ _00084_ _00002_ VGND VGND VPWR VPWR _00179_ sky130_fd_sc_hd__and2b_1
XFILLER_0_43_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_536 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08066_ _00108_ _00109_ VGND VGND VPWR VPWR _00110_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07729__B1 _06820_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13711__A1_N _02427_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08968_ _01072_ _01078_ VGND VGND VPWR VPWR _01079_ sky130_fd_sc_hd__xor2_1
X_07919_ _07046_ _07047_ net60 net3 VGND VGND VPWR VPWR _07048_ sky130_fd_sc_hd__and4bb_1
X_08899_ _01002_ _01003_ VGND VGND VPWR VPWR _01004_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10930_ _02520_ _03226_ _03228_ VGND VGND VPWR VPWR _03229_ sky130_fd_sc_hd__nor3_1
X_10861_ _03141_ _03144_ VGND VGND VPWR VPWR _03153_ sky130_fd_sc_hd__xor2_1
XFILLER_0_39_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12600_ _05061_ _05064_ VGND VGND VPWR VPWR _05065_ sky130_fd_sc_hd__or2b_1
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13580_ _01414_ _03783_ _06124_ VGND VGND VPWR VPWR _06125_ sky130_fd_sc_hd__and3_1
X_10792_ _05588_ _01933_ _03075_ _03076_ VGND VGND VPWR VPWR _03077_ sky130_fd_sc_hd__and4_1
XFILLER_0_109_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07530__A _04598_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13251__B _05773_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12531_ _04982_ _04987_ _04932_ VGND VGND VPWR VPWR _04989_ sky130_fd_sc_hd__a21oi_1
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10594__C _02856_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12462_ _04907_ _04912_ VGND VGND VPWR VPWR _04913_ sky130_fd_sc_hd__xnor2_2
XANTENNA__12005__A2 _02090_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07680__A2 net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_398 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14201_ _00344_ _00410_ VGND VGND VPWR VPWR _06793_ sky130_fd_sc_hd__nand2_2
X_11413_ _00268_ _01178_ _01248_ _06733_ VGND VGND VPWR VPWR _03759_ sky130_fd_sc_hd__a22o_1
X_12393_ _04834_ _04836_ VGND VGND VPWR VPWR _04837_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11764__A1 _02135_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14132_ _06657_ _06717_ _06716_ _06722_ VGND VGND VPWR VPWR _06729_ sky130_fd_sc_hd__a31o_1
XFILLER_0_105_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11344_ _03682_ VGND VGND VPWR VPWR _03683_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__08361__A _00414_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14063_ _06096_ _06653_ _06651_ VGND VGND VPWR VPWR _06655_ sky130_fd_sc_hd__nor3_1
X_11275_ _03604_ _03607_ VGND VGND VPWR VPWR _03608_ sky130_fd_sc_hd__and2_1
X_13014_ _05493_ _05494_ VGND VGND VPWR VPWR _05520_ sky130_fd_sc_hd__nand2_1
X_10226_ _02454_ _02455_ VGND VGND VPWR VPWR _02457_ sky130_fd_sc_hd__nand2_1
X_10157_ _02184_ _02208_ _02380_ VGND VGND VPWR VPWR _02381_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12611__A _00389_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10088_ _02304_ VGND VGND VPWR VPWR _02305_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_89_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13916_ _06361_ _06311_ _06359_ VGND VGND VPWR VPWR _06495_ sky130_fd_sc_hd__nor3_1
XANTENNA__10131__A _00151_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09893__B1 _02088_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09920__A _01361_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07143__C net61 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13847_ _02189_ _03783_ _05370_ VGND VGND VPWR VPWR _06419_ sky130_fd_sc_hd__and3_1
XFILLER_0_69_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13778_ _06335_ _06338_ _06341_ _06342_ VGND VGND VPWR VPWR _06343_ sky130_fd_sc_hd__a211o_1
XANTENNA__13441__A1 _01250_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08536__A _00605_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13441__B2 _01182_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07440__A net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13799__D _03683_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12729_ _05193_ _05195_ VGND VGND VPWR VPWR _05207_ sky130_fd_sc_hd__or2_1
XANTENNA__11452__B1 _02134_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08255__B _00159_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11897__A _06417_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap134 _06504_ VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__clkbuf_1
Xmax_cap145 _00313_ VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__clkbuf_1
XANTENNA__12505__B _03773_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09940_ _02111_ _02141_ VGND VGND VPWR VPWR _02143_ sky130_fd_sc_hd__and2_1
XFILLER_0_111_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12224__C _01248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09871_ _02063_ _02066_ VGND VGND VPWR VPWR _02067_ sky130_fd_sc_hd__xor2_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10025__B _02235_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08822_ _01044_ _05731_ net8 net9 VGND VGND VPWR VPWR _00919_ sky130_fd_sc_hd__and4_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13336__B _00745_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12878__D _02117_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08753_ _00670_ VGND VGND VPWR VPWR _00844_ sky130_fd_sc_hd__buf_4
XFILLER_0_24_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07704_ _01230_ _00475_ _06832_ VGND VGND VPWR VPWR _06833_ sky130_fd_sc_hd__and3_1
XTAP_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08684_ _00639_ _04015_ _04103_ _00563_ VGND VGND VPWR VPWR _00768_ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07635_ _06296_ _06307_ VGND VGND VPWR VPWR _06318_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_800 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07566_ _02664_ VGND VGND VPWR VPWR _05577_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_48_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09305_ _01329_ _01343_ VGND VGND VPWR VPWR _01447_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07497_ _04730_ _04796_ _04807_ VGND VGND VPWR VPWR _04818_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_63_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09236_ _01370_ _01371_ VGND VGND VPWR VPWR _01373_ sky130_fd_sc_hd__or2_1
XFILLER_0_134_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09167_ _01294_ _01296_ VGND VGND VPWR VPWR _01297_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09277__A _00431_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08118_ _00061_ _00161_ VGND VGND VPWR VPWR _00162_ sky130_fd_sc_hd__xor2_1
XFILLER_0_32_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08611__A1 _06428_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__08611__B2 _06450_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09098_ _01204_ _01220_ VGND VGND VPWR VPWR _01222_ sky130_fd_sc_hd__and2_1
XANTENNA__11957__D _03681_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08612__C _00144_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08049_ _00091_ _00092_ VGND VGND VPWR VPWR _00093_ sky130_fd_sc_hd__or2b_1
XFILLER_0_102_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11060_ _03278_ _03288_ VGND VGND VPWR VPWR _03372_ sky130_fd_sc_hd__and2_1
XANTENNA__07178__A1 _01284_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10011_ _01709_ _01881_ _01880_ VGND VGND VPWR VPWR _02221_ sky130_fd_sc_hd__a21o_1
XANTENNA__07178__B2 _01230_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11962_ _03059_ _03678_ _04361_ VGND VGND VPWR VPWR _04363_ sky130_fd_sc_hd__a21oi_1
XANTENNA__13671__A1 _01183_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09162__D _01288_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10485__A1 _02247_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13701_ _02426_ _02721_ _06246_ VGND VGND VPWR VPWR _06258_ sky130_fd_sc_hd__a21oi_1
X_10913_ _02534_ _03160_ VGND VGND VPWR VPWR _03210_ sky130_fd_sc_hd__and2_1
XFILLER_0_98_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10485__B2 _01473_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11893_ _04255_ _04286_ VGND VGND VPWR VPWR _04287_ sky130_fd_sc_hd__xnor2_2
X_13632_ _06048_ _06073_ VGND VGND VPWR VPWR _06182_ sky130_fd_sc_hd__nand2_1
X_10844_ _03129_ _03131_ _03133_ VGND VGND VPWR VPWR _03134_ sky130_fd_sc_hd__o21a_1
XFILLER_0_67_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13563_ _06074_ _04014_ _06104_ _06105_ VGND VGND VPWR VPWR _06106_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_137_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10775_ _03056_ _03057_ VGND VGND VPWR VPWR _03058_ sky130_fd_sc_hd__xnor2_1
X_12514_ _04968_ _04969_ VGND VGND VPWR VPWR _04970_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_137_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13494_ _06028_ _06029_ VGND VGND VPWR VPWR _06030_ sky130_fd_sc_hd__nand2_1
XANTENNA__08850__A1 _02664_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07653__A2 _06472_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07410__D _03718_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12445_ _04892_ _04891_ VGND VGND VPWR VPWR _04894_ sky130_fd_sc_hd__and2b_1
XFILLER_0_34_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07405__A2 _03685_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12376_ _04801_ _04806_ VGND VGND VPWR VPWR _04819_ sky130_fd_sc_hd__xnor2_1
X_14115_ _06700_ _06710_ VGND VGND VPWR VPWR _06711_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10771__D _02727_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08522__C _03707_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07810__C1 _06938_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11327_ _03638_ _03665_ VGND VGND VPWR VPWR _03666_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14046_ _06594_ _06592_ VGND VGND VPWR VPWR _06638_ sky130_fd_sc_hd__nor2_1
XANTENNA_output76_A net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11258_ _03577_ _03589_ _03575_ VGND VGND VPWR VPWR _03590_ sky130_fd_sc_hd__o21ba_1
X_10209_ _02424_ _02437_ VGND VGND VPWR VPWR _02438_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09634__B _04510_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11189_ _03508_ _03513_ _03509_ _03506_ VGND VGND VPWR VPWR _03514_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_89_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07420_ _03916_ _03960_ VGND VGND VPWR VPWR _03971_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_427 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07892__A2 _03499_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07170__A net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07351_ _03125_ _03191_ VGND VGND VPWR VPWR _03213_ sky130_fd_sc_hd__and2_4
XFILLER_0_128_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12219__C _01180_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07282_ _02335_ VGND VGND VPWR VPWR _02456_ sky130_fd_sc_hd__buf_4
XFILLER_0_17_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09021_ _06964_ _06966_ _00142_ _04895_ VGND VGND VPWR VPWR _01137_ sky130_fd_sc_hd__and4_1
XFILLER_0_127_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12235__B _00778_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10036__A _00844_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10951__A2 _01508_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09825__A _03510_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09923_ _02114_ _02123_ VGND VGND VPWR VPWR _02124_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09854_ _02047_ _01633_ _02048_ VGND VGND VPWR VPWR _02049_ sky130_fd_sc_hd__a21oi_4
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11900__A1 _02040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07345__A net61 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08805_ _03850_ _04510_ net13 _00730_ VGND VGND VPWR VPWR _00900_ sky130_fd_sc_hd__and4_1
XANTENNA__11900__B2 _02135_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09785_ _01961_ _01962_ _01971_ VGND VGND VPWR VPWR _01973_ sky130_fd_sc_hd__or3_1
X_08736_ _00377_ _00114_ _06765_ _02993_ VGND VGND VPWR VPWR _00826_ sky130_fd_sc_hd__a22o_1
XTAP_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08667_ _00587_ _00588_ _00749_ VGND VGND VPWR VPWR _00750_ sky130_fd_sc_hd__o21bai_2
XTAP_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07618_ _06065_ _06076_ _06120_ VGND VGND VPWR VPWR _06131_ sky130_fd_sc_hd__nand3b_4
XTAP_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12208__A2 _01954_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13513__C _02736_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08598_ _00669_ _00674_ VGND VGND VPWR VPWR _00675_ sky130_fd_sc_hd__xor2_1
XFILLER_0_49_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07549_ _04961_ _05379_ VGND VGND VPWR VPWR _05390_ sky130_fd_sc_hd__xnor2_2
XANTENNA__09085__A1 _02127_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10560_ _00294_ _01934_ VGND VGND VPWR VPWR _02822_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09219_ _01310_ _01352_ VGND VGND VPWR VPWR _01354_ sky130_fd_sc_hd__or2b_1
XFILLER_0_106_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10491_ _02741_ _02745_ VGND VGND VPWR VPWR _02746_ sky130_fd_sc_hd__xor2_2
XFILLER_0_133_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12230_ _01517_ _03748_ _04657_ VGND VGND VPWR VPWR _04658_ sky130_fd_sc_hd__and3_1
XFILLER_0_32_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_675 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12161_ _04473_ _04483_ VGND VGND VPWR VPWR _04582_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08060__A2 _00101_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11112_ _03423_ _03427_ _03428_ VGND VGND VPWR VPWR _03429_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_102_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09735__A _01339_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12092_ _04432_ _04504_ VGND VGND VPWR VPWR _04506_ sky130_fd_sc_hd__nor2_1
X_11043_ _02569_ _02572_ _03352_ VGND VGND VPWR VPWR _03353_ sky130_fd_sc_hd__a21o_1
XANTENNA__07255__A _02149_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12994_ _05497_ _05022_ _00381_ _02008_ VGND VGND VPWR VPWR _05498_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_87_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11945_ _04342_ _04343_ VGND VGND VPWR VPWR _04344_ sky130_fd_sc_hd__and2_1
XFILLER_0_86_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07702__B net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11876_ _04256_ _04267_ VGND VGND VPWR VPWR _04269_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13615_ _06152_ _06162_ VGND VGND VPWR VPWR _06163_ sky130_fd_sc_hd__and2b_1
XANTENNA__11407__B1 _03748_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10827_ _03111_ _03115_ VGND VGND VPWR VPWR _03116_ sky130_fd_sc_hd__nor2_1
XFILLER_0_144_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13546_ _06085_ _06086_ VGND VGND VPWR VPWR _06088_ sky130_fd_sc_hd__xor2_1
XFILLER_0_137_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07626__A2 _00650_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10758_ _03023_ _03039_ VGND VGND VPWR VPWR _03040_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08823__A1 _01044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08823__B2 _05731_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13477_ _06009_ _01956_ _03687_ _01414_ VGND VGND VPWR VPWR _06012_ sky130_fd_sc_hd__a22o_1
XFILLER_0_124_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10689_ _05203_ _01058_ _02962_ _02963_ VGND VGND VPWR VPWR _02964_ sky130_fd_sc_hd__a31o_1
XFILLER_0_35_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12428_ _04827_ _04875_ VGND VGND VPWR VPWR _04876_ sky130_fd_sc_hd__or2_1
XFILLER_0_113_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12359_ _00742_ _00605_ VGND VGND VPWR VPWR _04800_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14029_ _06618_ _06580_ VGND VGND VPWR VPWR _06619_ sky130_fd_sc_hd__xor2_2
X_09570_ _01456_ _01463_ VGND VGND VPWR VPWR _01738_ sky130_fd_sc_hd__nand2_1
X_08521_ _03059_ _00389_ _00393_ _02280_ VGND VGND VPWR VPWR _00590_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08708__B net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11415__A _06775_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08452_ _00514_ _00512_ VGND VGND VPWR VPWR _00515_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07403_ _00322_ _03773_ VGND VGND VPWR VPWR _03784_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08383_ _00417_ _00438_ VGND VGND VPWR VPWR _00439_ sky130_fd_sc_hd__xor2_4
XFILLER_0_58_594 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07334_ _02138_ _00410_ _03015_ _00333_ VGND VGND VPWR VPWR _03026_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_91_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09539__B _02960_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07265_ _02259_ _00333_ VGND VGND VPWR VPWR _02270_ sky130_fd_sc_hd__and2_2
XFILLER_0_61_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12246__A _04037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09004_ _01020_ _01023_ _01007_ VGND VGND VPWR VPWR _01118_ sky130_fd_sc_hd__o21a_1
XFILLER_0_116_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07196_ _00420_ _00978_ _00705_ _01208_ VGND VGND VPWR VPWR _01514_ sky130_fd_sc_hd__and4_1
XFILLER_0_5_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09906_ _02103_ _02104_ VGND VGND VPWR VPWR _02106_ sky130_fd_sc_hd__nand2_1
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09837_ _01980_ _02030_ VGND VGND VPWR VPWR _02031_ sky130_fd_sc_hd__xnor2_2
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09768_ _01954_ VGND VGND VPWR VPWR _01955_ sky130_fd_sc_hd__buf_4
XANTENNA__07526__A2_N _04378_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08719_ _03532_ _00121_ _04895_ _04873_ VGND VGND VPWR VPWR _00807_ sky130_fd_sc_hd__and4_1
XTAP_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09699_ _01872_ _01878_ VGND VGND VPWR VPWR _01879_ sky130_fd_sc_hd__xor2_1
XFILLER_0_69_848 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07522__B net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11730_ _04107_ _04057_ VGND VGND VPWR VPWR _04108_ sky130_fd_sc_hd__nor2_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10586__D _02304_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11661_ _04029_ _04031_ VGND VGND VPWR VPWR _04032_ sky130_fd_sc_hd__nand2_1
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13400_ _05913_ _05927_ VGND VGND VPWR VPWR _05928_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10612_ _02852_ _02847_ VGND VGND VPWR VPWR _02879_ sky130_fd_sc_hd__or2b_1
XFILLER_0_119_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11592_ _03955_ VGND VGND VPWR VPWR _03956_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_789 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13331_ _05411_ _05415_ VGND VGND VPWR VPWR _05852_ sky130_fd_sc_hd__or2b_1
XFILLER_0_52_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10543_ _00388_ _03004_ _02724_ _02727_ VGND VGND VPWR VPWR _02803_ sky130_fd_sc_hd__and4_1
XFILLER_0_91_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13262_ _05778_ _05786_ VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__xnor2_4
X_10474_ net57 VGND VGND VPWR VPWR _02727_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_121_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12213_ _00605_ _01507_ _01179_ _01254_ VGND VGND VPWR VPWR _04639_ sky130_fd_sc_hd__and4_1
XFILLER_0_121_135 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13193_ _05716_ VGND VGND VPWR VPWR _05717_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12144_ _00530_ _01183_ VGND VGND VPWR VPWR _04563_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12075_ _04452_ _04453_ VGND VGND VPWR VPWR _04487_ sky130_fd_sc_hd__nor2_1
XANTENNA__10404__A _02007_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10679__A1 _02982_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11026_ _03313_ _03315_ _03333_ _03309_ VGND VGND VPWR VPWR _03335_ sky130_fd_sc_hd__a211o_1
XANTENNA__11219__B _01108_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10679__B2 _00377_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07713__A _00880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12977_ _03602_ _05479_ VGND VGND VPWR VPWR _05480_ sky130_fd_sc_hd__xor2_2
XANTENNA__11880__D _00916_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10777__C _02723_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11928_ _03932_ _04325_ VGND VGND VPWR VPWR _04326_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10496__D _02731_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11859_ _04234_ _04243_ VGND VGND VPWR VPWR _04250_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08544__A _01372_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13529_ _06066_ _06067_ VGND VGND VPWR VPWR _06069_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput103 net103 VGND VGND VPWR VPWR prod[44] sky130_fd_sc_hd__clkbuf_4
Xoutput114 net114 VGND VGND VPWR VPWR prod[54] sky130_fd_sc_hd__clkbuf_4
Xoutput125 net125 VGND VGND VPWR VPWR prod[6] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_140_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_656 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12513__B _00755_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07952_ _07079_ _07080_ VGND VGND VPWR VPWR _07081_ sky130_fd_sc_hd__xor2_2
XANTENNA__11867__B1 _00575_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07883_ net177 net149 net39 net38 VGND VGND VPWR VPWR _07012_ sky130_fd_sc_hd__and4_1
X_09622_ _01791_ _01794_ VGND VGND VPWR VPWR _01795_ sky130_fd_sc_hd__xor2_1
XANTENNA__09822__B net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08719__A _03532_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10968__B net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09553_ _01482_ VGND VGND VPWR VPWR _01719_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08438__B _05478_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08504_ net14 VGND VGND VPWR VPWR _00571_ sky130_fd_sc_hd__buf_2
X_09484_ _01641_ _01432_ _01642_ VGND VGND VPWR VPWR _01643_ sky130_fd_sc_hd__o21ai_2
XANTENNA__12292__B1 _02189_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08435_ _00172_ _00174_ _00324_ _00495_ VGND VGND VPWR VPWR _00496_ sky130_fd_sc_hd__a31o_2
XFILLER_0_77_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_851 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08366_ _02127_ _03894_ _03872_ _03861_ VGND VGND VPWR VPWR _00421_ sky130_fd_sc_hd__a31o_1
X_07317_ _01853_ _02489_ _02828_ VGND VGND VPWR VPWR _02839_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_33_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08297_ _00252_ _00253_ _00343_ VGND VGND VPWR VPWR _00346_ sky130_fd_sc_hd__nor3_1
XFILLER_0_18_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08263__A2 _00143_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12407__C _00413_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07248_ _01569_ net181 VGND VGND VPWR VPWR _02083_ sky130_fd_sc_hd__xor2_2
XFILLER_0_61_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08015__A2 net6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07179_ _01262_ _01273_ _01317_ VGND VGND VPWR VPWR _01328_ sky130_fd_sc_hd__and3_1
XANTENNA__11030__D _00613_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10358__B1 _00423_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10190_ _02415_ _02416_ VGND VGND VPWR VPWR _02417_ sky130_fd_sc_hd__or2_1
XANTENNA__07517__B _05027_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12900_ _05230_ _05393_ VGND VGND VPWR VPWR _05395_ sky130_fd_sc_hd__nand2_1
XANTENNA__13535__A _01958_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13880_ _06438_ _06441_ VGND VGND VPWR VPWR _06455_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07533__A _01405_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12796__D _02723_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12831_ _05307_ _05310_ VGND VGND VPWR VPWR _05319_ sky130_fd_sc_hd__nand2_1
XTAP_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12762_ _04645_ _04646_ _05242_ VGND VGND VPWR VPWR _05243_ sky130_fd_sc_hd__nor3_1
XTAP_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11713_ _04084_ _04085_ _04088_ VGND VGND VPWR VPWR _04089_ sky130_fd_sc_hd__o21a_1
XFILLER_0_68_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12693_ _04694_ _05166_ VGND VGND VPWR VPWR _05167_ sky130_fd_sc_hd__nor2_1
XTAP_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13270__A _05779_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11644_ _03699_ VGND VGND VPWR VPWR _04013_ sky130_fd_sc_hd__buf_2
XFILLER_0_83_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput16 a[23] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__dlymetal6s2s_1
X_11575_ _00263_ _03750_ VGND VGND VPWR VPWR _03937_ sky130_fd_sc_hd__nand2_1
Xinput27 a[4] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13420__D _01250_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput38 b[14] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__buf_4
XFILLER_0_80_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13314_ _05679_ _05694_ _05712_ VGND VGND VPWR VPWR _05835_ sky130_fd_sc_hd__nand3_1
XFILLER_0_91_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08514__D _03938_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10526_ _02782_ _02783_ VGND VGND VPWR VPWR _02785_ sky130_fd_sc_hd__nand2_1
Xinput49 b[24] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10118__B _02190_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13245_ _05548_ _05557_ _05560_ VGND VGND VPWR VPWR _05770_ sky130_fd_sc_hd__and3_1
X_10457_ _02704_ _02705_ _02707_ VGND VGND VPWR VPWR _02710_ sky130_fd_sc_hd__nand3_1
XFILLER_0_32_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08811__B net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07708__A net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13176_ _05479_ _04608_ _04611_ _05697_ _04621_ VGND VGND VPWR VPWR _05699_ sky130_fd_sc_hd__o311a_1
X_10388_ _02617_ _02633_ VGND VGND VPWR VPWR _02634_ sky130_fd_sc_hd__xor2_1
X_12127_ _04541_ _04544_ VGND VGND VPWR VPWR _04545_ sky130_fd_sc_hd__and2_1
X_12058_ _04458_ _04465_ _04468_ VGND VGND VPWR VPWR _04469_ sky130_fd_sc_hd__o21ba_1
XANTENNA__13445__A _01183_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11009_ _05203_ _00604_ _02549_ _02548_ _01369_ VGND VGND VPWR VPWR _03316_ sky130_fd_sc_hd__a32o_1
XANTENNA__08539__A _00453_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12274__B1 _03686_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08220_ _06472_ _06483_ _00262_ _00263_ VGND VGND VPWR VPWR _00264_ sky130_fd_sc_hd__and4_1
XFILLER_0_56_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_564 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08705__C net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08151_ net150 _06175_ _06406_ VGND VGND VPWR VPWR _00195_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11412__B _06765_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09442__A1 _06439_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09442__B2 _02018_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07102_ _00475_ VGND VGND VPWR VPWR _00486_ sky130_fd_sc_hd__clkbuf_4
X_08082_ _00124_ _00125_ VGND VGND VPWR VPWR _00126_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_31_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09817__B _02008_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08984_ _00954_ _01094_ VGND VGND VPWR VPWR _01096_ sky130_fd_sc_hd__and2_1
X_07935_ _07058_ _07063_ VGND VGND VPWR VPWR _07064_ sky130_fd_sc_hd__xor2_1
X_07866_ _06991_ _06992_ _06994_ VGND VGND VPWR VPWR _06995_ sky130_fd_sc_hd__a21oi_1
X_09605_ _01774_ _01775_ VGND VGND VPWR VPWR _01776_ sky130_fd_sc_hd__or2_1
X_07797_ _06923_ _06924_ _06925_ VGND VGND VPWR VPWR _06926_ sky130_fd_sc_hd__or3_4
X_09536_ _01698_ _01699_ VGND VGND VPWR VPWR _01701_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07503__D _04873_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09467_ _01307_ _01625_ VGND VGND VPWR VPWR _01626_ sky130_fd_sc_hd__xor2_4
XFILLER_0_65_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08418_ _06472_ _00003_ _00270_ _00269_ VGND VGND VPWR VPWR _00478_ sky130_fd_sc_hd__a31o_1
XFILLER_0_93_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_862 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09398_ _01372_ net49 VGND VGND VPWR VPWR _01550_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12418__B _00378_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08349_ _00186_ _00402_ VGND VGND VPWR VPWR _00403_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_123_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_191 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11360_ _03695_ _03692_ _03698_ _03700_ VGND VGND VPWR VPWR _03701_ sky130_fd_sc_hd__nor4_1
XANTENNA__09984__A2 _02188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10311_ _02971_ _01368_ _00959_ _00366_ VGND VGND VPWR VPWR _02549_ sky130_fd_sc_hd__a22o_1
X_11291_ _03456_ _03496_ _03625_ VGND VGND VPWR VPWR _03626_ sky130_fd_sc_hd__or3_2
XFILLER_0_30_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13030_ _04603_ _05537_ VGND VGND VPWR VPWR _05538_ sky130_fd_sc_hd__xor2_2
X_10242_ _02086_ _02108_ _02144_ VGND VGND VPWR VPWR _02474_ sky130_fd_sc_hd__a21bo_1
XANTENNA__11695__D _01211_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10173_ _02069_ _02071_ _02068_ VGND VGND VPWR VPWR _02398_ sky130_fd_sc_hd__a21o_1
XFILLER_0_28_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13932_ _06481_ _06451_ _06479_ VGND VGND VPWR VPWR _06512_ sky130_fd_sc_hd__nor3_1
XANTENNA__08359__A net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13863_ _06434_ _06435_ VGND VGND VPWR VPWR _06436_ sky130_fd_sc_hd__nor2_1
XANTENNA__13048__A2 _00391_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10401__B _05467_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08078__B _00121_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12814_ _05090_ _05117_ VGND VGND VPWR VPWR _05300_ sky130_fd_sc_hd__and2_1
XANTENNA__08509__D _00571_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13794_ _06289_ _06262_ _06287_ VGND VGND VPWR VPWR _06360_ sky130_fd_sc_hd__nor3_1
XFILLER_0_69_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12745_ _05222_ _05223_ VGND VGND VPWR VPWR _05224_ sky130_fd_sc_hd__xor2_1
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12609__A _00915_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08094__A _05478_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12676_ _00381_ _01958_ _05146_ _04718_ VGND VGND VPWR VPWR _05149_ sky130_fd_sc_hd__a211o_1
XFILLER_0_25_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12328__B _01188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11627_ _03958_ _03968_ VGND VGND VPWR VPWR _03995_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11232__B _03559_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_139 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09918__A _02117_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11558_ _03897_ _03918_ VGND VGND VPWR VPWR _03919_ sky130_fd_sc_hd__or2_1
XFILLER_0_40_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08822__A _01044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10509_ _02765_ VGND VGND VPWR VPWR _02766_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__09637__B net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11489_ _03840_ _03842_ VGND VGND VPWR VPWR _03843_ sky130_fd_sc_hd__and2b_1
XFILLER_0_0_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09188__B1 _00294_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07438__A _00978_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13228_ _05528_ _05582_ _05586_ VGND VGND VPWR VPWR _05755_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_21_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07157__B net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13159_ _05648_ _05679_ VGND VGND VPWR VPWR _05680_ sky130_fd_sc_hd__nand2_1
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10742__B1 _01414_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09075__D net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07720_ _06841_ _06847_ _06848_ VGND VGND VPWR VPWR _06849_ sky130_fd_sc_hd__a21o_1
X_07651_ _06483_ VGND VGND VPWR VPWR _06494_ sky130_fd_sc_hd__buf_4
X_07582_ _05731_ _01000_ _00628_ _05742_ VGND VGND VPWR VPWR _05753_ sky130_fd_sc_hd__and4_1
X_09321_ _01447_ _01464_ VGND VGND VPWR VPWR _01465_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08466__A2 _00095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09252_ _01388_ _01389_ VGND VGND VPWR VPWR _01390_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12238__B _02120_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08203_ _06998_ _00203_ VGND VGND VPWR VPWR _00247_ sky130_fd_sc_hd__and2_1
XFILLER_0_44_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11142__B _03449_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09183_ _01312_ _00543_ _00636_ _00526_ VGND VGND VPWR VPWR _01314_ sky130_fd_sc_hd__and4_1
XFILLER_0_28_394 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_448 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08134_ _00100_ _00177_ VGND VGND VPWR VPWR _00178_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08732__A _00262_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07977__A1 _02719_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08065_ _00006_ _00107_ VGND VGND VPWR VPWR _00109_ sky130_fd_sc_hd__or2_1
XFILLER_0_70_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09547__B _01712_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07729__A1 net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07729__B2 _00563_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08967_ _01075_ _01077_ VGND VGND VPWR VPWR _01078_ sky130_fd_sc_hd__xnor2_2
X_07918_ net62 net61 net32 net2 VGND VGND VPWR VPWR _07047_ sky130_fd_sc_hd__and4_1
XANTENNA__12486__B1 _00741_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10502__A _01934_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08898_ _00997_ _01001_ VGND VGND VPWR VPWR _01003_ sky130_fd_sc_hd__or2_1
X_07849_ _06856_ _06882_ VGND VGND VPWR VPWR _06978_ sky130_fd_sc_hd__nand2_1
X_10860_ _03150_ _03151_ VGND VGND VPWR VPWR _03152_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_78_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09519_ _01502_ _01510_ _01512_ _01371_ VGND VGND VPWR VPWR _01682_ sky130_fd_sc_hd__a211oi_2
XANTENNA__07811__A net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10791_ _02149_ net54 _02312_ _02105_ VGND VGND VPWR VPWR _03076_ sky130_fd_sc_hd__a22o_1
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12530_ _04932_ _04982_ _04987_ VGND VGND VPWR VPWR _04988_ sky130_fd_sc_hd__and3_1
XFILLER_0_94_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10594__D _02858_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12461_ _04908_ _04911_ VGND VGND VPWR VPWR _04912_ sky130_fd_sc_hd__nor2_1
XFILLER_0_124_506 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_139 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14200_ _02401_ _06792_ VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__nor2_2
X_11412_ _00114_ _06765_ _01179_ _01254_ VGND VGND VPWR VPWR _03758_ sky130_fd_sc_hd__nand4_1
XFILLER_0_50_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12392_ _01517_ _01780_ _04835_ VGND VGND VPWR VPWR _04836_ sky130_fd_sc_hd__and3_1
X_14131_ _06699_ _06728_ VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__xor2_4
XFILLER_0_22_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11343_ _03681_ VGND VGND VPWR VPWR _03682_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_120_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14062_ _06096_ _06651_ _06653_ VGND VGND VPWR VPWR _06654_ sky130_fd_sc_hd__o21a_1
X_11274_ _03606_ VGND VGND VPWR VPWR _03607_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13013_ _05509_ _05517_ _05518_ VGND VGND VPWR VPWR _05519_ sky130_fd_sc_hd__o21a_2
X_10225_ _02113_ _02453_ VGND VGND VPWR VPWR _02455_ sky130_fd_sc_hd__nand2_1
X_10156_ _02184_ _02208_ _02235_ VGND VGND VPWR VPWR _02380_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_146_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12611__B _00393_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10087_ _02156_ VGND VGND VPWR VPWR _02304_ sky130_fd_sc_hd__buf_2
XFILLER_0_55_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13915_ _06488_ _06490_ VGND VGND VPWR VPWR _06493_ sky130_fd_sc_hd__nor2_1
XANTENNA__10131__B _01517_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09893__A1 _06626_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09893__B2 _06450_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09920__B _00159_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13846_ _05902_ _05905_ VGND VGND VPWR VPWR _06418_ sky130_fd_sc_hd__nor2_1
XANTENNA__07143__D net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08817__A _00742_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13442__B _02765_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13777_ _06339_ _06327_ VGND VGND VPWR VPWR _06342_ sky130_fd_sc_hd__nor2_1
X_10989_ _03260_ _03293_ VGND VGND VPWR VPWR _03294_ sky130_fd_sc_hd__nand2_1
XANTENNA__12339__A _00755_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13441__A2 _02721_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11452__A1 _06964_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12728_ _05202_ _05205_ VGND VGND VPWR VPWR _05206_ sky130_fd_sc_hd__or2_4
XANTENNA__11452__B2 _06966_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__08255__C _00144_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12659_ _05118_ _05129_ VGND VGND VPWR VPWR _05130_ sky130_fd_sc_hd__xor2_2
XFILLER_0_127_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11897__B _06439_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap135 _06583_ VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__buf_1
Xmax_cap146 _04265_ VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__clkbuf_1
XANTENNA__09086__C _00730_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09870_ _02064_ _02065_ VGND VGND VPWR VPWR _02066_ sky130_fd_sc_hd__nand2_1
XANTENNA__12224__D _02117_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09383__A _06472_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08821_ _00747_ _00750_ VGND VGND VPWR VPWR _00918_ sky130_fd_sc_hd__and2_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08752_ _00257_ VGND VGND VPWR VPWR _00843_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__13336__C _02724_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07703_ net149 net63 _06830_ _06831_ VGND VGND VPWR VPWR _06832_ sky130_fd_sc_hd__a31o_1
X_08683_ _00563_ _00639_ _04015_ _04103_ VGND VGND VPWR VPWR _00767_ sky130_fd_sc_hd__and4_1
X_07634_ _05868_ _05901_ _06285_ VGND VGND VPWR VPWR _06307_ sky130_fd_sc_hd__and3_1
XFILLER_0_17_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08483__B1_N _00342_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07565_ _03268_ VGND VGND VPWR VPWR _05566_ sky130_fd_sc_hd__buf_4
XANTENNA__09636__A1 _01177_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_812 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09304_ _01311_ _01352_ VGND VGND VPWR VPWR _01446_ sky130_fd_sc_hd__and2b_1
XFILLER_0_36_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07496_ _04642_ _04708_ _04719_ VGND VGND VPWR VPWR _04807_ sky130_fd_sc_hd__o21a_1
XFILLER_0_61_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09235_ _01284_ _01230_ _01368_ _00959_ VGND VGND VPWR VPWR _01371_ sky130_fd_sc_hd__and4_1
XFILLER_0_106_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09166_ _01189_ _01225_ _01224_ VGND VGND VPWR VPWR _01296_ sky130_fd_sc_hd__a21o_1
XFILLER_0_44_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08462__A _07040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08117_ _00157_ _00158_ _00160_ VGND VGND VPWR VPWR _00161_ sky130_fd_sc_hd__and3_1
XFILLER_0_121_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09277__B _04169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09097_ _01204_ _01220_ VGND VGND VPWR VPWR _01221_ sky130_fd_sc_hd__nor2_1
XANTENNA__08611__A2 _00144_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08048_ _03521_ _02993_ _06875_ _00377_ VGND VGND VPWR VPWR _00092_ sky130_fd_sc_hd__a22o_1
XANTENNA__08612__D _00298_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07178__A2 _01295_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10010_ _02218_ _02219_ VGND VGND VPWR VPWR _02220_ sky130_fd_sc_hd__and2b_1
X_09999_ _02206_ _02207_ VGND VGND VPWR VPWR _02208_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_98_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11961_ _03059_ _03678_ _04361_ VGND VGND VPWR VPWR _04362_ sky130_fd_sc_hd__and3_1
XANTENNA__13671__A2 _02766_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10912_ _03131_ _03208_ VGND VGND VPWR VPWR _03209_ sky130_fd_sc_hd__nor2_1
X_13700_ _06254_ _06256_ VGND VGND VPWR VPWR _06257_ sky130_fd_sc_hd__nor2_1
XANTENNA__10485__A2 _02736_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11892_ _04284_ _04285_ VGND VGND VPWR VPWR _04286_ sky130_fd_sc_hd__nor2_1
XANTENNA__08637__A _00598_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13631_ _06048_ _06073_ VGND VGND VPWR VPWR _06181_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10843_ _03124_ _03132_ VGND VGND VPWR VPWR _03133_ sky130_fd_sc_hd__nor2_1
XANTENNA__13262__B _05786_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13562_ _06075_ _06077_ _06078_ _02736_ VGND VGND VPWR VPWR _06105_ sky130_fd_sc_hd__nand4_1
X_10774_ _06494_ _02168_ VGND VGND VPWR VPWR _03057_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12513_ _04059_ _00755_ VGND VGND VPWR VPWR _04969_ sky130_fd_sc_hd__nand2_2
XFILLER_0_81_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13493_ _06024_ _06027_ VGND VGND VPWR VPWR _06029_ sky130_fd_sc_hd__or2_1
XFILLER_0_82_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08850__A2 net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12444_ _04891_ _04892_ VGND VGND VPWR VPWR _04893_ sky130_fd_sc_hd__and2b_1
XFILLER_0_35_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12375_ _04815_ _04816_ VGND VGND VPWR VPWR _04817_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10407__A _02029_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14114_ _06708_ _06709_ VGND VGND VPWR VPWR _06710_ sky130_fd_sc_hd__and2_1
XFILLER_0_50_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08522__D _00392_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11326_ _03640_ _03663_ VGND VGND VPWR VPWR _03665_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14045_ _06533_ _06596_ VGND VGND VPWR VPWR _06636_ sky130_fd_sc_hd__xnor2_2
X_11257_ _03580_ _03545_ _03581_ VGND VGND VPWR VPWR _03589_ sky130_fd_sc_hd__nand3_1
XFILLER_0_66_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08366__A1 _02127_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10208_ _02433_ _02436_ VGND VGND VPWR VPWR _02437_ sky130_fd_sc_hd__xnor2_2
XANTENNA_output69_A net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11188_ net138 _03505_ VGND VGND VPWR VPWR _03513_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09634__C net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12341__B _03762_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10139_ _00457_ _02224_ _02360_ VGND VGND VPWR VPWR _02361_ sky130_fd_sc_hd__and3_1
XANTENNA__09931__A net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13453__A _03783_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13829_ _06397_ _06398_ VGND VGND VPWR VPWR _06399_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07350_ _03125_ _03191_ VGND VGND VPWR VPWR _03202_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07281_ _01985_ _02423_ _02434_ VGND VGND VPWR VPWR _02445_ sky130_fd_sc_hd__a21o_1
XANTENNA__12219__D _01249_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09020_ _06966_ _00142_ VGND VGND VPWR VPWR _01136_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12235__C _01178_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09922_ _02115_ _02122_ VGND VGND VPWR VPWR _02123_ sky130_fd_sc_hd__xor2_1
XANTENNA__09825__B net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09853_ _01833_ _01834_ VGND VGND VPWR VPWR _02048_ sky130_fd_sc_hd__nand2_1
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11900__A2 _03681_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08804_ _00889_ _00892_ VGND VGND VPWR VPWR _00899_ sky130_fd_sc_hd__or2b_4
X_09784_ _01961_ _01962_ _01971_ VGND VGND VPWR VPWR _01972_ sky130_fd_sc_hd__o21a_1
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_92 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08735_ _00822_ _00823_ VGND VGND VPWR VPWR _00824_ sky130_fd_sc_hd__xnor2_1
XTAP_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13363__A _00416_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08666_ _00421_ _00427_ _00586_ VGND VGND VPWR VPWR _00749_ sky130_fd_sc_hd__and3_1
XANTENNA__11664__A1 _00575_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07617_ _06098_ _06109_ VGND VGND VPWR VPWR _06120_ sky130_fd_sc_hd__xor2_4
XTAP_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08597_ _00671_ _00673_ VGND VGND VPWR VPWR _00674_ sky130_fd_sc_hd__nor2_1
XTAP_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09609__A1 _02040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09609__B2 _00415_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13513__D _02737_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07548_ _04972_ _04840_ VGND VGND VPWR VPWR _05379_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09085__A2 _00734_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07479_ net162 net44 net31 net32 VGND VGND VPWR VPWR _04620_ sky130_fd_sc_hd__and4_1
XFILLER_0_64_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09218_ _01311_ _01352_ VGND VGND VPWR VPWR _01353_ sky130_fd_sc_hd__xor2_1
XFILLER_0_134_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10490_ _02247_ _02742_ _02744_ VGND VGND VPWR VPWR _02745_ sky130_fd_sc_hd__and3_1
XFILLER_0_44_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09149_ _01274_ _01275_ _01209_ _01212_ VGND VGND VPWR VPWR _01277_ sky130_fd_sc_hd__a211oi_1
X_12160_ _04471_ _04485_ VGND VGND VPWR VPWR _04581_ sky130_fd_sc_hd__nor2_4
XFILLER_0_114_391 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11111_ _02561_ _03424_ _03426_ VGND VGND VPWR VPWR _03428_ sky130_fd_sc_hd__o21a_1
X_12091_ _04432_ _04504_ VGND VGND VPWR VPWR _04505_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11042_ _00158_ _04059_ _02570_ VGND VGND VPWR VPWR _03352_ sky130_fd_sc_hd__and3_1
XFILLER_0_36_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12993_ _05021_ VGND VGND VPWR VPWR _05497_ sky130_fd_sc_hd__inv_2
XANTENNA__12852__B1 _02305_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11944_ _04340_ _04341_ _04269_ VGND VGND VPWR VPWR _04343_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07271__A _02280_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07702__C net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11875_ net146 _04266_ VGND VGND VPWR VPWR _04267_ sky130_fd_sc_hd__nor2_1
X_13614_ _06152_ _06160_ _06161_ VGND VGND VPWR VPWR _06162_ sky130_fd_sc_hd__or3_1
X_10826_ _03112_ _03113_ VGND VGND VPWR VPWR _03115_ sky130_fd_sc_hd__or2_1
XANTENNA__11407__A1 _00257_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11407__B2 _00670_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13545_ _05985_ _02737_ _05995_ VGND VGND VPWR VPWR _06086_ sky130_fd_sc_hd__and3_1
X_10757_ _03024_ _03021_ VGND VGND VPWR VPWR _03039_ sky130_fd_sc_hd__or2_1
XANTENNA__08284__B1 _06875_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08823__A2 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13476_ _01414_ _06009_ _01956_ _03687_ VGND VGND VPWR VPWR _06011_ sky130_fd_sc_hd__and4_1
XFILLER_0_14_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10688_ _00366_ _02982_ net50 _01546_ VGND VGND VPWR VPWR _02963_ sky130_fd_sc_hd__and4_1
X_12427_ _04837_ _04872_ _04874_ VGND VGND VPWR VPWR _04875_ sky130_fd_sc_hd__o21ba_1
XANTENNA__10137__A _05203_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12358_ _04792_ _04791_ VGND VGND VPWR VPWR _04799_ sky130_fd_sc_hd__and2b_1
XFILLER_0_50_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11309_ _02913_ _03645_ VGND VGND VPWR VPWR _03646_ sky130_fd_sc_hd__nand2_1
XANTENNA__12352__A _03696_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12289_ _04707_ _04722_ VGND VGND VPWR VPWR _04723_ sky130_fd_sc_hd__xor2_1
X_14028_ _05417_ _05954_ _05955_ VGND VGND VPWR VPWR _06618_ sky130_fd_sc_hd__o21ai_2
XANTENNA__13167__B _05688_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10146__A1 _04851_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10146__B2 net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08520_ _00587_ net160 VGND VGND VPWR VPWR _00589_ sky130_fd_sc_hd__xor2_2
XANTENNA__10600__A _04862_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07181__A _01339_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08451_ _00296_ _00301_ VGND VGND VPWR VPWR _00514_ sky130_fd_sc_hd__and2_1
XFILLER_0_77_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11415__B _02119_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07402_ _03762_ VGND VGND VPWR VPWR _03773_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_86_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08382_ _00436_ _00437_ VGND VGND VPWR VPWR _00438_ sky130_fd_sc_hd__and2_1
XFILLER_0_45_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07333_ _03004_ VGND VGND VPWR VPWR _03015_ sky130_fd_sc_hd__buf_4
XFILLER_0_73_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_716 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07264_ _02116_ VGND VGND VPWR VPWR _02259_ sky130_fd_sc_hd__buf_4
XFILLER_0_116_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09539__C net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09003_ _01020_ _01023_ VGND VGND VPWR VPWR _01117_ sky130_fd_sc_hd__and2_1
XFILLER_0_61_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12246__B _00783_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07195_ _00420_ _01197_ _01208_ _00978_ VGND VGND VPWR VPWR _01503_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__08740__A _07004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xwire3 _06691_ VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__clkbuf_1
XANTENNA__14180__C _02742_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07356__A _02719_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09905_ _01995_ _02102_ VGND VGND VPWR VPWR _02104_ sky130_fd_sc_hd__nand2_1
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09836_ _02006_ _02028_ VGND VGND VPWR VPWR _02030_ sky130_fd_sc_hd__xor2_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09767_ _01953_ VGND VGND VPWR VPWR _01954_ sky130_fd_sc_hd__clkbuf_4
XTAP_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08718_ _00641_ _00805_ _00660_ VGND VGND VPWR VPWR _00806_ sky130_fd_sc_hd__a21oi_1
XTAP_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09698_ _01876_ _01877_ VGND VGND VPWR VPWR _01878_ sky130_fd_sc_hd__xnor2_1
XTAP_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07091__A _00355_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08649_ net14 VGND VGND VPWR VPWR _00730_ sky130_fd_sc_hd__buf_2
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07522__C _00355_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13821__A _04714_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11660_ _04006_ _04030_ VGND VGND VPWR VPWR _04031_ sky130_fd_sc_hd__xnor2_1
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10611_ _00310_ _01060_ _02869_ _02877_ VGND VGND VPWR VPWR _02878_ sky130_fd_sc_hd__a31o_1
X_11591_ _03891_ _03954_ VGND VGND VPWR VPWR _03955_ sky130_fd_sc_hd__xor2_1
XFILLER_0_52_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11341__A _03679_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_407 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13330_ _05318_ _05419_ VGND VGND VPWR VPWR _05851_ sky130_fd_sc_hd__and2b_1
X_10542_ _03004_ _02724_ _02728_ _00388_ VGND VGND VPWR VPWR _02802_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13261_ _02278_ _05756_ _05781_ _05782_ _05785_ VGND VGND VPWR VPWR _05786_ sky130_fd_sc_hd__a311o_4
XFILLER_0_134_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10473_ _02725_ VGND VGND VPWR VPWR _02726_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_106_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08569__A1 _03543_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12212_ _04636_ _04637_ VGND VGND VPWR VPWR _04638_ sky130_fd_sc_hd__xnor2_1
X_13192_ _05464_ _05466_ VGND VGND VPWR VPWR _05716_ sky130_fd_sc_hd__nand2_1
XANTENNA__08650__A _04510_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10376__A1 _00413_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12143_ _04558_ _04559_ _04561_ VGND VGND VPWR VPWR _04562_ sky130_fd_sc_hd__o21a_1
XFILLER_0_130_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__07266__A _02040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12074_ _04471_ _04484_ _04485_ VGND VGND VPWR VPWR _04486_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_47_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10404__B _02117_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11025_ _03321_ _03331_ _03332_ VGND VGND VPWR VPWR _03333_ sky130_fd_sc_hd__o21a_1
XANTENNA__08741__A1 _00543_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07713__B net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12976_ _04606_ _04607_ _05477_ _04614_ VGND VGND VPWR VPWR _05479_ sky130_fd_sc_hd__o211a_1
XFILLER_0_99_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10777__D _02727_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11927_ _03930_ _03931_ VGND VGND VPWR VPWR _04325_ sky130_fd_sc_hd__or2_1
XFILLER_0_87_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11858_ _04236_ _04248_ VGND VGND VPWR VPWR _04249_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_86_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08825__A _01996_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13450__B _02722_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10809_ _03062_ _03058_ VGND VGND VPWR VPWR _03096_ sky130_fd_sc_hd__or2b_1
XFILLER_0_138_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11789_ _03850_ _01394_ net22 net24 VGND VGND VPWR VPWR _04173_ sky130_fd_sc_hd__and4_1
XANTENNA__08544__B _04268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13528_ _06066_ _06067_ VGND VGND VPWR VPWR _06068_ sky130_fd_sc_hd__nor2_1
XFILLER_0_125_431 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07480__A1 net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13459_ _05978_ _05991_ VGND VGND VPWR VPWR _05992_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09757__B1 _01712_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput104 net104 VGND VGND VPWR VPWR prod[45] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_70_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput115 net115 VGND VGND VPWR VPWR prod[55] sky130_fd_sc_hd__buf_2
XFILLER_0_140_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput126 net126 VGND VGND VPWR VPWR prod[7] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07176__A _01197_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07951_ _06935_ _06982_ _06981_ VGND VGND VPWR VPWR _07080_ sky130_fd_sc_hd__a21boi_4
XFILLER_0_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07882_ _00978_ _07010_ net38 net149 VGND VGND VPWR VPWR _07011_ sky130_fd_sc_hd__a22oi_1
XANTENNA__11867__A1 _00113_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11867__B2 _00258_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09621_ _01792_ _01793_ VGND VGND VPWR VPWR _01794_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08719__B _00121_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09552_ _01716_ _01717_ VGND VGND VPWR VPWR _01718_ sky130_fd_sc_hd__xor2_1
XANTENNA__10968__C net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08503_ _00417_ _00436_ _00437_ VGND VGND VPWR VPWR _00570_ sky130_fd_sc_hd__a21bo_1
XANTENNA__08438__C _00142_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09483_ _01428_ _01431_ VGND VGND VPWR VPWR _01642_ sky130_fd_sc_hd__nand2_1
XANTENNA__08496__B1 _04004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12292__A1 _02187_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12292__B2 _00575_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08434_ _00325_ _00494_ _00323_ VGND VGND VPWR VPWR _00495_ sky130_fd_sc_hd__a21o_1
XFILLER_0_86_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08365_ _03916_ _03960_ VGND VGND VPWR VPWR _00419_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_705 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_280 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07316_ _02806_ _02817_ VGND VGND VPWR VPWR _02828_ sky130_fd_sc_hd__nor2_1
X_08296_ _00252_ _00253_ _00343_ VGND VGND VPWR VPWR _00345_ sky130_fd_sc_hd__o21a_1
XFILLER_0_61_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07247_ _01011_ _02061_ VGND VGND VPWR VPWR _02072_ sky130_fd_sc_hd__nor2_1
XANTENNA__12407__D _00571_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07178_ _01284_ _01295_ _01306_ _01230_ VGND VGND VPWR VPWR _01317_ sky130_fd_sc_hd__a22o_1
XANTENNA__08470__A _03532_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10358__A1 _07010_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10358__B2 _00101_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07086__A _00300_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07814__A _00541_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09819_ _01765_ _01769_ VGND VGND VPWR VPWR _02011_ sky130_fd_sc_hd__and2_1
XANTENNA__07533__B _05203_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12830_ _03676_ _05317_ _02792_ _04600_ VGND VGND VPWR VPWR _05318_ sky130_fd_sc_hd__a31o_1
XTAP_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12761_ _05238_ _05241_ VGND VGND VPWR VPWR _05242_ sky130_fd_sc_hd__xnor2_1
XTAP_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11712_ _04051_ _04087_ VGND VGND VPWR VPWR _04088_ sky130_fd_sc_hd__xor2_1
XTAP_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_487 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12692_ _04692_ _04693_ VGND VGND VPWR VPWR _05166_ sky130_fd_sc_hd__nor2_1
XANTENNA__08645__A _00725_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11643_ _03859_ _04009_ _04011_ VGND VGND VPWR VPWR _04012_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_127_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11574_ _03934_ _03935_ VGND VGND VPWR VPWR _03936_ sky130_fd_sc_hd__or2b_1
XFILLER_0_80_833 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput17 a[24] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_2
Xinput28 a[5] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__buf_6
XFILLER_0_91_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput39 b[15] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__buf_2
XANTENNA__07462__A1 net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10525_ _02774_ _02779_ _02781_ VGND VGND VPWR VPWR _02783_ sky130_fd_sc_hd__nand3_1
XFILLER_0_107_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13313_ _05663_ _05834_ VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__xnor2_2
XFILLER_0_52_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13244_ _02713_ _05579_ _05768_ VGND VGND VPWR VPWR _05769_ sky130_fd_sc_hd__and3_1
X_10456_ _02704_ _02705_ _02707_ VGND VGND VPWR VPWR _02709_ sky130_fd_sc_hd__a21o_2
XFILLER_0_110_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13175_ _03613_ _03623_ _04616_ VGND VGND VPWR VPWR _05697_ sky130_fd_sc_hd__nand3_1
XANTENNA__07708__B net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10387_ _02630_ _02632_ VGND VGND VPWR VPWR _02633_ sky130_fd_sc_hd__or2_1
X_12126_ _04001_ _04542_ VGND VGND VPWR VPWR _04544_ sky130_fd_sc_hd__and2_1
XANTENNA__08962__A1 _04081_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12057_ _04458_ _04465_ _04467_ VGND VGND VPWR VPWR _04468_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_74_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11008_ _00294_ _01505_ _03314_ VGND VGND VPWR VPWR _03315_ sky130_fd_sc_hd__and3_1
XFILLER_0_74_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13445__B _01252_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08539__B _02051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12274__A1 _00376_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12959_ _04536_ _04454_ VGND VGND VPWR VPWR _05460_ sky130_fd_sc_hd__nand2_1
XANTENNA__12274__B2 _00380_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_142_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10037__B1 _02247_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08150_ _05313_ _00193_ VGND VGND VPWR VPWR _00194_ sky130_fd_sc_hd__xor2_2
XANTENNA__08705__D net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11412__C _01179_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09089__C _01744_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09442__A2 _00414_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07101_ net63 VGND VGND VPWR VPWR _00475_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_15_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08081_ _00028_ _00030_ _00026_ VGND VGND VPWR VPWR _00125_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_141_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07205__A1 _01076_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08721__C _00497_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10325__A _04862_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08983_ _00954_ _01094_ VGND VGND VPWR VPWR _01095_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07934_ net172 _07062_ VGND VGND VPWR VPWR _07063_ sky130_fd_sc_hd__nor2_1
X_07865_ _06977_ _06993_ VGND VGND VPWR VPWR _06994_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08181__A2 _03609_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09604_ _06417_ _00138_ _00414_ _00574_ VGND VGND VPWR VPWR _01775_ sky130_fd_sc_hd__and4_1
X_07796_ _04532_ _05225_ _04499_ VGND VGND VPWR VPWR _06925_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_64_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09535_ _00355_ _02960_ _04180_ _04191_ VGND VGND VPWR VPWR _01699_ sky130_fd_sc_hd__and4_1
XANTENNA__10995__A _02247_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09466_ _01563_ _01623_ VGND VGND VPWR VPWR _01625_ sky130_fd_sc_hd__xor2_4
XFILLER_0_47_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08417_ _00474_ _00476_ VGND VGND VPWR VPWR _00477_ sky130_fd_sc_hd__xor2_1
X_09397_ _01546_ _01418_ _01548_ VGND VGND VPWR VPWR _01549_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_108_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12418__C _00414_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08348_ _06999_ _00363_ _00360_ _00362_ VGND VGND VPWR VPWR _00402_ sky130_fd_sc_hd__o22a_1
XFILLER_0_74_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_833 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08279_ _00172_ _00174_ _00325_ VGND VGND VPWR VPWR _00326_ sky130_fd_sc_hd__a21o_1
XFILLER_0_144_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10310_ _00366_ _02971_ _01368_ VGND VGND VPWR VPWR _02548_ sky130_fd_sc_hd__and3_1
XANTENNA__07809__A _06626_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11290_ _03536_ _03616_ _03621_ _03624_ _03495_ VGND VGND VPWR VPWR _03625_ sky130_fd_sc_hd__o311a_1
X_10241_ _02438_ _02472_ VGND VGND VPWR VPWR _02473_ sky130_fd_sc_hd__xnor2_1
X_10172_ _02395_ _02396_ VGND VGND VPWR VPWR _02397_ sky130_fd_sc_hd__nor2_1
XFILLER_0_100_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13480__A1_N _01108_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13931_ _06359_ _06510_ VGND VGND VPWR VPWR _06511_ sky130_fd_sc_hd__nor2_1
X_13862_ _06431_ _06432_ VGND VGND VPWR VPWR _06435_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12813_ _05295_ _05298_ VGND VGND VPWR VPWR _05299_ sky130_fd_sc_hd__xnor2_1
X_13793_ _06328_ _06356_ _06358_ VGND VGND VPWR VPWR _06359_ sky130_fd_sc_hd__o21a_1
XFILLER_0_139_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12744_ _00375_ _03681_ VGND VGND VPWR VPWR _05223_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12609__B _01059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12675_ _05146_ _04718_ _00381_ _01958_ VGND VGND VPWR VPWR _05147_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_65_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12328__C _03414_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11626_ _03984_ _03990_ _03992_ VGND VGND VPWR VPWR _03994_ sky130_fd_sc_hd__or3_1
XFILLER_0_37_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11557_ _03521_ _02117_ _03895_ _03896_ VGND VGND VPWR VPWR _03918_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_69_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08822__B _05731_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10508_ _02759_ VGND VGND VPWR VPWR _02765_ sky130_fd_sc_hd__clkbuf_4
X_11488_ _03722_ _03841_ VGND VGND VPWR VPWR _03842_ sky130_fd_sc_hd__and2_1
XFILLER_0_123_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_590 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09188__A1 _00257_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09188__B2 _00670_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10439_ _02688_ _02689_ VGND VGND VPWR VPWR _02690_ sky130_fd_sc_hd__or2_2
X_13227_ _05424_ _05754_ VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__xor2_1
XANTENNA__11773__A2_N _01960_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13158_ _05663_ _05678_ VGND VGND VPWR VPWR _05679_ sky130_fd_sc_hd__and2_4
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10742__B2 _07040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12109_ _04500_ _04502_ _04524_ VGND VGND VPWR VPWR _04525_ sky130_fd_sc_hd__a21oi_4
X_13089_ _05492_ _05597_ _05602_ VGND VGND VPWR VPWR _05603_ sky130_fd_sc_hd__a21bo_1
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07454__A _01996_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13692__B1 _02737_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07650_ _05566_ VGND VGND VPWR VPWR _06483_ sky130_fd_sc_hd__clkbuf_4
X_07581_ _00639_ VGND VGND VPWR VPWR _05742_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__12247__A1 _00378_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09112__A1 _00943_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09320_ _01456_ _01463_ VGND VGND VPWR VPWR _01464_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09251_ _01086_ _01092_ _01387_ VGND VGND VPWR VPWR _01389_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_8_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08202_ _00244_ _00239_ _00202_ VGND VGND VPWR VPWR _00246_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09182_ _00544_ _00636_ _00526_ _01312_ VGND VGND VPWR VPWR _01313_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08133_ _00081_ _00176_ VGND VGND VPWR VPWR _00177_ sky130_fd_sc_hd__xor2_1
XFILLER_0_71_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08732__B _00818_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07977__A2 _03499_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08064_ _00006_ _00107_ VGND VGND VPWR VPWR _00108_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07729__A2 net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08966_ _04268_ net46 VGND VGND VPWR VPWR _01077_ sky130_fd_sc_hd__nand2_1
X_07917_ net62 net32 _04367_ net61 VGND VGND VPWR VPWR _07046_ sky130_fd_sc_hd__a22oi_1
XANTENNA__12486__A1 _00779_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08897_ _00997_ _01001_ VGND VGND VPWR VPWR _01002_ sky130_fd_sc_hd__nand2_1
XANTENNA__12486__B2 _00783_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07848_ _06893_ VGND VGND VPWR VPWR _06977_ sky130_fd_sc_hd__inv_2
X_07779_ _06904_ _06907_ VGND VGND VPWR VPWR _06908_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09518_ _01515_ _01524_ VGND VGND VPWR VPWR _01681_ sky130_fd_sc_hd__nand2_1
XANTENNA__07811__B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10790_ _03074_ VGND VGND VPWR VPWR _03075_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_90 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09449_ _01292_ _01604_ VGND VGND VPWR VPWR _01606_ sky130_fd_sc_hd__and2_1
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_800 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12460_ _04903_ _04904_ VGND VGND VPWR VPWR _04911_ sky130_fd_sc_hd__and2_1
XFILLER_0_124_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11411_ _03747_ _03756_ VGND VGND VPWR VPWR _03757_ sky130_fd_sc_hd__or2b_1
XFILLER_0_124_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12391_ _01518_ _01601_ VGND VGND VPWR VPWR _04835_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14130_ _06726_ _06727_ VGND VGND VPWR VPWR _06728_ sky130_fd_sc_hd__nand2_2
X_11342_ _02459_ VGND VGND VPWR VPWR _03681_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__10972__A1 _00145_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14061_ _06085_ _06086_ _06090_ _06652_ VGND VGND VPWR VPWR _06653_ sky130_fd_sc_hd__a211o_1
X_11273_ _03572_ _03560_ _03605_ VGND VGND VPWR VPWR _03606_ sky130_fd_sc_hd__o21a_1
X_13012_ _05510_ _05516_ VGND VGND VPWR VPWR _05518_ sky130_fd_sc_hd__nand2_1
X_10224_ _02113_ _02453_ VGND VGND VPWR VPWR _02454_ sky130_fd_sc_hd__or2_1
X_10155_ _02347_ _02377_ VGND VGND VPWR VPWR _02378_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12611__C _01060_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10086_ _02155_ _02161_ VGND VGND VPWR VPWR _02303_ sky130_fd_sc_hd__and2_1
XFILLER_0_89_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13914_ _06240_ _06188_ _06491_ VGND VGND VPWR VPWR _06492_ sky130_fd_sc_hd__mux2_2
XANTENNA__09893__A2 _02090_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13845_ _06411_ _06415_ VGND VGND VPWR VPWR _06416_ sky130_fd_sc_hd__nor2_1
XANTENNA__09920__C _02119_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13776_ _06339_ _06326_ _06325_ VGND VGND VPWR VPWR _06341_ sky130_fd_sc_hd__o21a_1
X_10988_ _03259_ _03255_ VGND VGND VPWR VPWR _03293_ sky130_fd_sc_hd__or2b_1
XFILLER_0_146_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12339__B _01260_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12727_ _05191_ _05204_ VGND VGND VPWR VPWR _05205_ sky130_fd_sc_hd__xnor2_2
XANTENNA__11452__A2 _01953_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__08255__D _00298_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12658_ _05125_ _05128_ VGND VGND VPWR VPWR _05129_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11609_ _00654_ _01181_ _01250_ _00543_ VGND VGND VPWR VPWR _03975_ sky130_fd_sc_hd__a22o_1
XANTENNA__11897__C _01954_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12589_ _00745_ _01412_ _05044_ _05043_ VGND VGND VPWR VPWR _05053_ sky130_fd_sc_hd__a31o_1
XFILLER_0_111_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09086__D net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08908__A1 _06775_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08908__B2 _00258_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08820_ _00157_ _00159_ _00915_ _00916_ VGND VGND VPWR VPWR _00917_ sky130_fd_sc_hd__and4_1
XANTENNA__12090__A _06626_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09383__B _00458_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07184__A _01372_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08751_ _00686_ _00703_ VGND VGND VPWR VPWR _00842_ sky130_fd_sc_hd__nand2_1
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13336__D _02728_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07702_ net1 net12 net64 net34 VGND VGND VPWR VPWR _06831_ sky130_fd_sc_hd__and4_1
X_08682_ _00603_ _00624_ _00625_ VGND VGND VPWR VPWR _00766_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_136_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07912__A _02456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07633_ _05868_ _05901_ _06285_ VGND VGND VPWR VPWR _06296_ sky130_fd_sc_hd__a21oi_1
X_07564_ _03279_ _03290_ _03301_ VGND VGND VPWR VPWR _05555_ sky130_fd_sc_hd__and3_1
XFILLER_0_88_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09303_ _01348_ _01351_ VGND VGND VPWR VPWR _01445_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_824 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_243 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07495_ _04774_ _04785_ VGND VGND VPWR VPWR _04796_ sky130_fd_sc_hd__and2_2
XFILLER_0_0_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09234_ _04268_ _01368_ _01369_ _01372_ VGND VGND VPWR VPWR _01370_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_134_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09165_ _01287_ _01293_ VGND VGND VPWR VPWR _01294_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08116_ _00159_ _00142_ VGND VGND VPWR VPWR _00160_ sky130_fd_sc_hd__nand2_1
XANTENNA__07359__A _01295_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09096_ _01217_ _01218_ VGND VGND VPWR VPWR _01220_ sky130_fd_sc_hd__nand2_1
XANTENNA__09277__C net50 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08047_ _03521_ _00377_ _02982_ _06875_ VGND VGND VPWR VPWR _00091_ sky130_fd_sc_hd__and4_1
XFILLER_0_4_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09998_ _01912_ _01915_ _01910_ VGND VGND VPWR VPWR _02207_ sky130_fd_sc_hd__a21o_1
XANTENNA__07583__B1 _05742_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07094__A _00388_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08949_ net49 VGND VGND VPWR VPWR _01058_ sky130_fd_sc_hd__buf_2
XFILLER_0_98_313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11960_ _04358_ _04360_ VGND VGND VPWR VPWR _04361_ sky130_fd_sc_hd__nor2_1
X_10911_ _02517_ _03130_ VGND VGND VPWR VPWR _03208_ sky130_fd_sc_hd__and2_1
X_11891_ _04102_ _04283_ _04282_ VGND VGND VPWR VPWR _04285_ sky130_fd_sc_hd__o21a_1
XFILLER_0_67_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11344__A _03682_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13630_ _06177_ _06179_ VGND VGND VPWR VPWR _06180_ sky130_fd_sc_hd__or2_1
XANTENNA__07541__B _05291_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10842_ _03119_ _03122_ _03123_ VGND VGND VPWR VPWR _03132_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_67_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13561_ _06077_ _06078_ _02736_ _01958_ VGND VGND VPWR VPWR _06104_ sky130_fd_sc_hd__a22o_1
X_10773_ _03054_ _03055_ VGND VGND VPWR VPWR _03056_ sky130_fd_sc_hd__or2b_1
XFILLER_0_54_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12512_ _04956_ _04955_ VGND VGND VPWR VPWR _04968_ sky130_fd_sc_hd__or2b_2
XFILLER_0_137_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09749__A _01933_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13492_ _06024_ _06027_ VGND VGND VPWR VPWR _06028_ sky130_fd_sc_hd__nand2_1
XANTENNA__08653__A net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12443_ _04876_ _04877_ VGND VGND VPWR VPWR _04892_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_136_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12374_ _00389_ _00392_ _00457_ _00607_ VGND VGND VPWR VPWR _04816_ sky130_fd_sc_hd__and4_1
XANTENNA__10407__B _01960_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14113_ _06663_ _06665_ _06707_ VGND VGND VPWR VPWR _06709_ sky130_fd_sc_hd__or3_1
XFILLER_0_120_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11325_ _03654_ _03662_ _03651_ VGND VGND VPWR VPWR _03663_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_22_379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11256_ _02299_ _02241_ _02384_ _03586_ _03584_ VGND VGND VPWR VPWR _03588_ sky130_fd_sc_hd__a2111o_1
X_14044_ _06587_ _06634_ VGND VGND VPWR VPWR _06635_ sky130_fd_sc_hd__or2_2
XFILLER_0_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09563__A1 _00544_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08366__A2 _03894_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10207_ _02003_ _02005_ _02103_ _02435_ VGND VGND VPWR VPWR _02436_ sky130_fd_sc_hd__a31oi_4
X_11187_ _03498_ _03511_ VGND VGND VPWR VPWR _03512_ sky130_fd_sc_hd__and2_1
XFILLER_0_66_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12341__C _01368_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10138_ _02358_ _02359_ VGND VGND VPWR VPWR _02360_ sky130_fd_sc_hd__xor2_1
XANTENNA__13734__A _00915_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10069_ _02253_ _02283_ VGND VGND VPWR VPWR _02284_ sky130_fd_sc_hd__and2_1
XFILLER_0_82_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08828__A _00901_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13828_ _04714_ _03680_ _06396_ VGND VGND VPWR VPWR _06398_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13759_ _06309_ _06321_ VGND VGND VPWR VPWR _06322_ sky130_fd_sc_hd__or2_1
XFILLER_0_73_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07280_ _01886_ _01930_ _01963_ VGND VGND VPWR VPWR _02434_ sky130_fd_sc_hd__and3_1
XFILLER_0_127_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12235__D _01248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09394__A net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09921_ _02118_ _02121_ VGND VGND VPWR VPWR _02122_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09852_ _01627_ _01628_ _01629_ _01630_ VGND VGND VPWR VPWR _02047_ sky130_fd_sc_hd__o211ai_1
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08803_ _00893_ _00897_ _00894_ _00721_ VGND VGND VPWR VPWR _00898_ sky130_fd_sc_hd__o2bb2a_4
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09783_ _01964_ _01970_ VGND VGND VPWR VPWR _01971_ sky130_fd_sc_hd__xor2_1
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08734_ _00649_ _00652_ _00648_ VGND VGND VPWR VPWR _00823_ sky130_fd_sc_hd__o21bai_1
XANTENNA__08738__A _06885_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13363__B _01288_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08665_ _00744_ _00746_ VGND VGND VPWR VPWR _00747_ sky130_fd_sc_hd__and2b_1
XFILLER_0_49_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07616_ _03114_ _03411_ _03400_ VGND VGND VPWR VPWR _06109_ sky130_fd_sc_hd__a21o_1
XTAP_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08596_ _06472_ _06483_ _00113_ _00258_ VGND VGND VPWR VPWR _00673_ sky130_fd_sc_hd__and4_1
XFILLER_0_95_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09609__A2 _01600_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07547_ _05313_ _05346_ _05357_ VGND VGND VPWR VPWR _05368_ sky130_fd_sc_hd__o21ai_2
XANTENNA__13810__B1 _03686_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_805 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07478_ net163 net31 net32 net44 VGND VGND VPWR VPWR _04609_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09490__B1 net52 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09217_ _01348_ _01351_ VGND VGND VPWR VPWR _01352_ sky130_fd_sc_hd__xor2_2
XANTENNA__10508__A _02759_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07089__A _00333_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09148_ _01209_ _01212_ _01274_ _01275_ VGND VGND VPWR VPWR _01276_ sky130_fd_sc_hd__o211a_1
XFILLER_0_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09079_ _01192_ _01200_ VGND VGND VPWR VPWR _01201_ sky130_fd_sc_hd__xor2_1
XFILLER_0_31_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11110_ _02561_ _03424_ _03426_ VGND VGND VPWR VPWR _03427_ sky130_fd_sc_hd__nor3_1
X_12090_ _06626_ _03680_ _04359_ VGND VGND VPWR VPWR _04504_ sky130_fd_sc_hd__and3_1
XANTENNA__07817__A _02719_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11041_ _03346_ _03349_ _03350_ VGND VGND VPWR VPWR _03351_ sky130_fd_sc_hd__and3_1
XANTENNA__11339__A _02673_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11557__A2_N _02117_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12992_ _05493_ _05494_ _05495_ VGND VGND VPWR VPWR _05496_ sky130_fd_sc_hd__a21o_1
XFILLER_0_99_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11943_ _04340_ _04269_ _04341_ VGND VGND VPWR VPWR _04342_ sky130_fd_sc_hd__or3_1
XFILLER_0_87_828 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12852__A1 _01586_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12852__B2 _00574_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08367__B _04510_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11874_ _04260_ _04263_ _04264_ _04262_ VGND VGND VPWR VPWR _04266_ sky130_fd_sc_hd__o22a_1
XANTENNA__07702__D net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13613_ _06147_ net141 _06151_ VGND VGND VPWR VPWR _06161_ sky130_fd_sc_hd__nor3_1
X_10825_ _01339_ _02312_ net57 _04081_ VGND VGND VPWR VPWR _03113_ sky130_fd_sc_hd__a22oi_1
XANTENNA__11407__A2 _03750_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13544_ _06049_ _06050_ _06051_ VGND VGND VPWR VPWR _06085_ sky130_fd_sc_hd__and3_1
XANTENNA__08284__A1 _00377_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_142 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10756_ _03034_ _03036_ VGND VGND VPWR VPWR _03038_ sky130_fd_sc_hd__nand2_1
XANTENNA__08284__B2 _02993_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13475_ _02856_ VGND VGND VPWR VPWR _06009_ sky130_fd_sc_hd__buf_2
XFILLER_0_82_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10687_ _02982_ net50 _02158_ _00366_ VGND VGND VPWR VPWR _02962_ sky130_fd_sc_hd__a22o_1
XANTENNA__10418__A _01295_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12426_ _04834_ _04836_ _04832_ VGND VGND VPWR VPWR _04874_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_23_633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10137__B net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12357_ _04794_ _04797_ VGND VGND VPWR VPWR _04798_ sky130_fd_sc_hd__and2_1
XFILLER_0_77_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output81_A net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11308_ _03634_ _03644_ VGND VGND VPWR VPWR _03645_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12288_ _04709_ _04705_ VGND VGND VPWR VPWR _04722_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11249__A _03566_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14027_ _05839_ _06614_ _06616_ VGND VGND VPWR VPWR _06617_ sky130_fd_sc_hd__a21oi_2
X_11239_ _02980_ _03568_ VGND VGND VPWR VPWR _03569_ sky130_fd_sc_hd__nand2_1
XANTENNA__10146__A2 _04015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13464__A _01252_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13183__B _05688_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10600__B _04873_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08450_ _00296_ _00301_ _00512_ VGND VGND VPWR VPWR _00513_ sky130_fd_sc_hd__and3_2
XFILLER_0_89_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07401_ net10 VGND VGND VPWR VPWR _03762_ sky130_fd_sc_hd__clkbuf_4
X_08381_ _00434_ _00435_ VGND VGND VPWR VPWR _00437_ sky130_fd_sc_hd__or2_1
XFILLER_0_147_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07332_ _02993_ VGND VGND VPWR VPWR _03004_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_85_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10082__A1 _00991_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07263_ _02215_ _02237_ VGND VGND VPWR VPWR _02248_ sky130_fd_sc_hd__or2_1
XFILLER_0_116_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10328__A _05027_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09002_ _01027_ _01030_ VGND VGND VPWR VPWR _01116_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12246__C _01178_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07194_ _01459_ _01481_ VGND VGND VPWR VPWR _01492_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_130_104 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11031__B1 _00778_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_159 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09904_ _01995_ _02102_ VGND VGND VPWR VPWR _02103_ sky130_fd_sc_hd__or2_1
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09835_ _02009_ _02027_ VGND VGND VPWR VPWR _02028_ sky130_fd_sc_hd__xnor2_2
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09766_ net21 VGND VGND VPWR VPWR _01953_ sky130_fd_sc_hd__buf_2
X_08717_ _00653_ _00658_ VGND VGND VPWR VPWR _00805_ sky130_fd_sc_hd__or2b_1
XTAP_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09697_ _04598_ _04026_ VGND VGND VPWR VPWR _01877_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer40 _03246_ VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__dlygate4sd1_1
XTAP_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08648_ _00589_ _00590_ _00591_ _00728_ VGND VGND VPWR VPWR _00729_ sky130_fd_sc_hd__a31o_2
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07522__D _02960_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13821__B _03683_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08579_ _00004_ VGND VGND VPWR VPWR _00654_ sky130_fd_sc_hd__buf_4
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10610_ _02876_ VGND VGND VPWR VPWR _02877_ sky130_fd_sc_hd__inv_2
XANTENNA__08266__A1 _02280_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11590_ _03951_ _03953_ VGND VGND VPWR VPWR _03954_ sky130_fd_sc_hd__or2_2
XFILLER_0_9_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10541_ _02799_ _02800_ VGND VGND VPWR VPWR _02801_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13260_ _05772_ _05779_ _05784_ VGND VGND VPWR VPWR _05785_ sky130_fd_sc_hd__a21o_1
X_10472_ _02724_ VGND VGND VPWR VPWR _02725_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_32_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08569__A2 _00294_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12211_ _00376_ _00379_ _01954_ _02135_ VGND VGND VPWR VPWR _04637_ sky130_fd_sc_hd__and4_1
X_13191_ _05708_ _05714_ VGND VGND VPWR VPWR _05715_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_103_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08650__B _00661_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12142_ _04478_ _04560_ VGND VGND VPWR VPWR _04561_ sky130_fd_sc_hd__or2_1
XANTENNA__13268__B _05792_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12073_ _04457_ _04470_ VGND VGND VPWR VPWR _04485_ sky130_fd_sc_hd__nor2_1
X_11024_ _03313_ _03315_ VGND VGND VPWR VPWR _03332_ sky130_fd_sc_hd__xor2_1
XANTENNA__10701__A _00095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07282__A _02335_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12975_ _04602_ _04607_ VGND VGND VPWR VPWR _05477_ sky130_fd_sc_hd__or2_1
XFILLER_0_63_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11926_ _04253_ _04322_ VGND VGND VPWR VPWR _04324_ sky130_fd_sc_hd__nand2_1
XANTENNA__07701__B1 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11857_ _04242_ _04241_ VGND VGND VPWR VPWR _04248_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08825__B _03762_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10808_ _06494_ _01934_ _03086_ _03094_ VGND VGND VPWR VPWR _03095_ sky130_fd_sc_hd__a31o_1
XFILLER_0_55_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11788_ _02127_ net24 _02668_ _02667_ net21 VGND VGND VPWR VPWR _04172_ sky130_fd_sc_hd__a32o_1
XFILLER_0_82_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08544__C _00612_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13527_ _06031_ _06046_ _06044_ VGND VGND VPWR VPWR _06067_ sky130_fd_sc_hd__a21oi_1
X_10739_ _02986_ _02973_ _02984_ VGND VGND VPWR VPWR _03019_ sky130_fd_sc_hd__and3_1
XFILLER_0_137_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13458_ _05989_ _05990_ VGND VGND VPWR VPWR _05991_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07480__A2 _04367_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12409_ _04059_ _01584_ VGND VGND VPWR VPWR _04855_ sky130_fd_sc_hd__nand2_1
Xoutput105 net105 VGND VGND VPWR VPWR prod[46] sky130_fd_sc_hd__clkbuf_4
X_13389_ _00375_ _02673_ _05388_ _05387_ VGND VGND VPWR VPWR _05916_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_23_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput116 net116 VGND VGND VPWR VPWR prod[56] sky130_fd_sc_hd__buf_4
XFILLER_0_50_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput127 net127 VGND VGND VPWR VPWR prod[8] sky130_fd_sc_hd__clkbuf_4
XANTENNA__07457__A _04367_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07950_ _07077_ _07078_ VGND VGND VPWR VPWR _07079_ sky130_fd_sc_hd__nor2_1
X_07881_ net39 VGND VGND VPWR VPWR _07010_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__11867__A2 _00415_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09620_ _01275_ _01588_ _01592_ VGND VGND VPWR VPWR _01793_ sky130_fd_sc_hd__and3_1
XANTENNA__09415__A1_N _00322_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07192__A _00661_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09551_ _01360_ _01422_ _01557_ _01556_ _01493_ VGND VGND VPWR VPWR _01717_ sky130_fd_sc_hd__a32o_1
XANTENNA__10968__D _01368_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08719__C _04895_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08502_ _00567_ _00569_ VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__xnor2_4
X_09482_ _01243_ VGND VGND VPWR VPWR _01641_ sky130_fd_sc_hd__inv_2
XANTENNA__08438__D _04862_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12292__A2 _01601_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08433_ _00319_ _00320_ VGND VGND VPWR VPWR _00494_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08364_ _03949_ _03927_ VGND VGND VPWR VPWR _00418_ sky130_fd_sc_hd__or2b_1
XFILLER_0_129_771 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07315_ _02631_ _02795_ VGND VGND VPWR VPWR _02817_ sky130_fd_sc_hd__and2_1
XFILLER_0_34_717 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08295_ _00329_ _00342_ VGND VGND VPWR VPWR _00343_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_116_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09847__A _01828_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07246_ _00442_ _02018_ _02040_ _02051_ VGND VGND VPWR VPWR _02061_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_131_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_761 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11004__B1 _01369_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07177_ _01208_ VGND VGND VPWR VPWR _01306_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__08470__B _00151_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10358__A2 _03685_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11555__A1 _00486_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_833 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09818_ _00486_ _01260_ _01767_ VGND VGND VPWR VPWR _02010_ sky130_fd_sc_hd__and3_1
XANTENNA__07814__B _03499_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09749_ _01933_ VGND VGND VPWR VPWR _01934_ sky130_fd_sc_hd__clkbuf_4
XTAP_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12760_ _05239_ _05240_ VGND VGND VPWR VPWR _05241_ sky130_fd_sc_hd__xnor2_1
XTAP_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ _00257_ _00916_ _04086_ VGND VGND VPWR VPWR _04087_ sky130_fd_sc_hd__and3_1
XTAP_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12691_ _05162_ _05164_ VGND VGND VPWR VPWR _05165_ sky130_fd_sc_hd__xnor2_2
XTAP_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11352__A _01155_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11642_ _03844_ _04010_ VGND VGND VPWR VPWR _04011_ sky130_fd_sc_hd__and2_1
XTAP_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11573_ _03904_ _03911_ VGND VGND VPWR VPWR _03935_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput18 a[25] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_80_845 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13312_ _05830_ _05833_ VGND VGND VPWR VPWR _05834_ sky130_fd_sc_hd__nor2_1
XFILLER_0_134_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10524_ _02774_ _02779_ _02781_ VGND VGND VPWR VPWR _02782_ sky130_fd_sc_hd__a21o_1
Xinput29 a[6] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__buf_4
XFILLER_0_135_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08661__A _00159_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13243_ _05573_ _05767_ _05562_ VGND VGND VPWR VPWR _05768_ sky130_fd_sc_hd__and3b_2
X_10455_ _02389_ _02706_ _02388_ VGND VGND VPWR VPWR _02707_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_33_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11546__A1 _03532_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08411__A1 _06494_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13174_ _05691_ _05695_ VGND VGND VPWR VPWR _05696_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_0_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10386_ _02418_ _02629_ VGND VGND VPWR VPWR _02632_ sky130_fd_sc_hd__and2_1
X_12125_ _04000_ _03969_ _03997_ VGND VGND VPWR VPWR _04542_ sky130_fd_sc_hd__or3_1
XANTENNA__08962__A2 _00604_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12056_ _03928_ _03929_ VGND VGND VPWR VPWR _04467_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10106__A1_N _05588_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11007_ _00293_ _01664_ VGND VGND VPWR VPWR _03314_ sky130_fd_sc_hd__nand2_1
XANTENNA__13445__C _02766_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08539__C _00458_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13742__A _02088_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12958_ _04589_ _04487_ _05458_ VGND VGND VPWR VPWR _05459_ sky130_fd_sc_hd__o21a_1
XFILLER_0_99_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12274__A2 _01955_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11909_ _04303_ _04304_ VGND VGND VPWR VPWR _04305_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12889_ _05224_ _05381_ _05382_ VGND VGND VPWR VPWR _05383_ sky130_fd_sc_hd__a21o_1
XTAP_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10037__A1 _02246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10037__B2 _02249_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11412__D _01254_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09089__D _01211_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07100_ _00453_ VGND VGND VPWR VPWR _00464_ sky130_fd_sc_hd__buf_4
X_08080_ _00120_ _00123_ VGND VGND VPWR VPWR _00124_ sky130_fd_sc_hd__xor2_2
XANTENNA__09667__A _00654_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08571__A _06965_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13601__A1_N _01414_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11537__A1 _06873_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11537__B2 _06874_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07187__A _01383_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07205__A2 net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08721__D _00142_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10325__B net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08982_ _01085_ _01093_ VGND VGND VPWR VPWR _01094_ sky130_fd_sc_hd__xor2_1
X_07933_ _01470_ net7 _07059_ _07060_ VGND VGND VPWR VPWR _07062_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__11437__A _00844_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07864_ _06890_ _06892_ VGND VGND VPWR VPWR _06993_ sky130_fd_sc_hd__nand2_1
X_09603_ _06428_ _00415_ _00574_ _06439_ VGND VGND VPWR VPWR _01774_ sky130_fd_sc_hd__a22oi_1
X_07795_ _05236_ _05258_ VGND VGND VPWR VPWR _06924_ sky130_fd_sc_hd__and2b_1
XFILLER_0_64_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09534_ _02971_ _04103_ _00777_ _00366_ VGND VGND VPWR VPWR _01698_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_64_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10995__B _02190_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07650__A _05566_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09465_ _01572_ _01622_ VGND VGND VPWR VPWR _01623_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_109_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08416_ _06483_ _00003_ VGND VGND VPWR VPWR _00476_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09396_ _04169_ net50 _01545_ _00431_ VGND VGND VPWR VPWR _01548_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08347_ _00344_ _00391_ VGND VGND VPWR VPWR _00401_ sky130_fd_sc_hd__and2_1
XANTENNA__12418__D _00572_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_845 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_558 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08278_ _00170_ _00171_ VGND VGND VPWR VPWR _00325_ sky130_fd_sc_hd__and2b_1
XFILLER_0_104_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07229_ _01853_ _01864_ VGND VGND VPWR VPWR _01875_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07809__B _06450_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07097__A _00420_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10240_ _02142_ _02471_ VGND VGND VPWR VPWR _02472_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_131_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13827__A _01066_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10171_ _02393_ _02394_ VGND VGND VPWR VPWR _02396_ sky130_fd_sc_hd__nor2_1
XANTENNA__11347__A _03686_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13930_ _06358_ _06328_ _06356_ VGND VGND VPWR VPWR _06510_ sky130_fd_sc_hd__nor3_1
X_13861_ _06431_ _06432_ VGND VGND VPWR VPWR _06434_ sky130_fd_sc_hd__and2_1
XANTENNA__11466__A1_N _03543_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12812_ _05297_ VGND VGND VPWR VPWR _05298_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13792_ _06311_ _06357_ VGND VGND VPWR VPWR _06358_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12743_ _01953_ _05220_ _05221_ VGND VGND VPWR VPWR _05222_ sky130_fd_sc_hd__a21bo_1
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12674_ _04717_ VGND VGND VPWR VPWR _05146_ sky130_fd_sc_hd__inv_2
XTAP_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11625_ _03979_ _03991_ VGND VGND VPWR VPWR _03992_ sky130_fd_sc_hd__xor2_2
XANTENNA__12328__D _01289_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11810__A _06439_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11556_ _00497_ _02120_ _03915_ VGND VGND VPWR VPWR _03917_ sky130_fd_sc_hd__and3_1
XANTENNA__08391__A _04268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__08822__C net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10507_ _01472_ _02759_ _02761_ _02763_ VGND VGND VPWR VPWR _02764_ sky130_fd_sc_hd__and4_1
XFILLER_0_80_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11487_ _03711_ _03712_ _03721_ VGND VGND VPWR VPWR _03841_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09188__A2 _00293_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13226_ _05604_ _05680_ _05713_ _05733_ _05752_ VGND VGND VPWR VPWR _05754_ sky130_fd_sc_hd__o41a_1
XFILLER_0_122_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10438_ _02684_ _02685_ _02683_ VGND VGND VPWR VPWR _02689_ sky130_fd_sc_hd__and3_1
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13157_ _05667_ _05677_ VGND VGND VPWR VPWR _05678_ sky130_fd_sc_hd__xor2_2
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10369_ _02407_ _02611_ VGND VGND VPWR VPWR _02613_ sky130_fd_sc_hd__and2_1
XANTENNA__12641__A _00916_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10742__A2 _01061_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12108_ _04409_ _04494_ _04497_ VGND VGND VPWR VPWR _04524_ sky130_fd_sc_hd__or3_1
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13088_ _05598_ _05600_ _05601_ VGND VGND VPWR VPWR _05602_ sky130_fd_sc_hd__a21o_1
X_12039_ _04427_ _04447_ VGND VGND VPWR VPWR _04448_ sky130_fd_sc_hd__xor2_2
XFILLER_0_18_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07454__B _00901_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13692__A1 _02426_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13692__B2 _02427_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07580_ _03147_ VGND VGND VPWR VPWR _05731_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__12247__A2 _02119_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09250_ _01086_ _01092_ _01387_ VGND VGND VPWR VPWR _01388_ sky130_fd_sc_hd__and3_1
XFILLER_0_75_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08201_ _00244_ _00239_ VGND VGND VPWR VPWR _00245_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_145_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09181_ _00654_ VGND VGND VPWR VPWR _01312_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_8_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08132_ _00137_ _00175_ VGND VGND VPWR VPWR _00176_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08063_ _00105_ _00106_ VGND VGND VPWR VPWR _00107_ sky130_fd_sc_hd__nor2_1
XFILLER_0_114_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07645__A _06417_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08965_ _01073_ _01074_ VGND VGND VPWR VPWR _01075_ sky130_fd_sc_hd__and2b_1
X_07916_ _01996_ _04378_ _06913_ _06912_ VGND VGND VPWR VPWR _07045_ sky130_fd_sc_hd__a31o_1
X_08896_ _00998_ _00999_ VGND VGND VPWR VPWR _01001_ sky130_fd_sc_hd__and2_1
XANTENNA__12486__A2 _00755_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10497__A1 _01473_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07847_ _06973_ _06975_ VGND VGND VPWR VPWR _06976_ sky130_fd_sc_hd__xnor2_1
X_07778_ _06905_ _06906_ VGND VGND VPWR VPWR _06907_ sky130_fd_sc_hd__xor2_1
XANTENNA__07380__A _03521_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09517_ _01677_ _01679_ VGND VGND VPWR VPWR _01680_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11446__B1 _03678_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07811__C _06818_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_116 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09448_ _01292_ _01604_ VGND VGND VPWR VPWR _01605_ sky130_fd_sc_hd__nor2_1
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_812 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09379_ _01527_ _01528_ VGND VGND VPWR VPWR _01529_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_171 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11410_ _03754_ _03755_ VGND VGND VPWR VPWR _03756_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12390_ _04831_ _04832_ _04833_ VGND VGND VPWR VPWR _04834_ sky130_fd_sc_hd__and3_1
XFILLER_0_117_593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11341_ _03679_ VGND VGND VPWR VPWR _03680_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_34_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10972__A2 _00460_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14060_ _05969_ _05985_ _02743_ _02742_ VGND VGND VPWR VPWR _06652_ sky130_fd_sc_hd__and4_1
XANTENNA__07586__A2_N _05588_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11272_ _03572_ _03560_ _03569_ VGND VGND VPWR VPWR _03605_ sky130_fd_sc_hd__a21o_1
X_13011_ _05510_ _05516_ VGND VGND VPWR VPWR _05517_ sky130_fd_sc_hd__nor2_1
X_10223_ _02451_ _02452_ VGND VGND VPWR VPWR _02453_ sky130_fd_sc_hd__or2_1
XANTENNA__10185__B1 _00730_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07555__A _05445_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10154_ _02233_ _02376_ VGND VGND VPWR VPWR _02377_ sky130_fd_sc_hd__xnor2_4
XANTENNA__12611__D _01412_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10085_ _02167_ _02170_ _02173_ _02300_ _02178_ VGND VGND VPWR VPWR _02301_ sky130_fd_sc_hd__a32o_1
XANTENNA__09770__A _01956_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13913_ _06488_ _06490_ VGND VGND VPWR VPWR _06491_ sky130_fd_sc_hd__and2_1
X_13844_ _06410_ _06409_ VGND VGND VPWR VPWR _06415_ sky130_fd_sc_hd__and2b_1
XANTENNA__09920__D _02120_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13775_ _06320_ _06322_ VGND VGND VPWR VPWR _06339_ sky130_fd_sc_hd__and2_1
X_10987_ _00310_ _00459_ _03283_ _03291_ VGND VGND VPWR VPWR _03292_ sky130_fd_sc_hd__a31o_1
XFILLER_0_139_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12339__C _01507_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12726_ _05186_ _05188_ VGND VGND VPWR VPWR _05204_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12657_ _05088_ _05127_ VGND VGND VPWR VPWR _05128_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_65_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11540__A _06819_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11608_ _03775_ VGND VGND VPWR VPWR _03974_ sky130_fd_sc_hd__inv_2
XFILLER_0_143_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12588_ _05047_ _05051_ VGND VGND VPWR VPWR _05052_ sky130_fd_sc_hd__or2b_1
XFILLER_0_142_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11897__D _02135_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_142_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11539_ _03895_ _03897_ VGND VGND VPWR VPWR _03898_ sky130_fd_sc_hd__nor2_1
XFILLER_0_111_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08369__B1 net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08908__A2 _00095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13209_ _05728_ _05730_ VGND VGND VPWR VPWR _05735_ sky130_fd_sc_hd__or2_1
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14189_ _06787_ _06620_ VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__xnor2_4
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07465__A _00661_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12090__B _03680_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08750_ _00839_ _00840_ VGND VGND VPWR VPWR _00841_ sky130_fd_sc_hd__and2_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07701_ net12 net64 net34 net1 VGND VGND VPWR VPWR _06830_ sky130_fd_sc_hd__a22o_1
X_08681_ _00596_ _00764_ VGND VGND VPWR VPWR _00765_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_136_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07344__A1 net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07632_ _06263_ _06274_ VGND VGND VPWR VPWR _06285_ sky130_fd_sc_hd__or2_1
XANTENNA__07912__B _07040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07563_ _03345_ _03367_ _03334_ VGND VGND VPWR VPWR _05544_ sky130_fd_sc_hd__a21oi_2
X_09302_ _01165_ _01353_ _01354_ VGND VGND VPWR VPWR _01444_ sky130_fd_sc_hd__o21a_1
XFILLER_0_75_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07494_ net154 net170 VGND VGND VPWR VPWR _04785_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_119_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_255 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09233_ _00959_ VGND VGND VPWR VPWR _01369_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_118_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_214 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09164_ _01290_ _01292_ VGND VGND VPWR VPWR _01293_ sky130_fd_sc_hd__and2_1
XFILLER_0_145_187 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08115_ _01405_ VGND VGND VPWR VPWR _00159_ sky130_fd_sc_hd__buf_4
XANTENNA__10403__A1 _01178_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10066__A _01752_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07359__B _01405_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09095_ _00910_ _01216_ VGND VGND VPWR VPWR _01218_ sky130_fd_sc_hd__or2_1
XFILLER_0_142_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08046_ _00087_ _00088_ _00086_ VGND VGND VPWR VPWR _00090_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_102_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_572 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09574__B _01741_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12281__A _01066_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11903__A1 _02335_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09997_ _02203_ _02205_ VGND VGND VPWR VPWR _02206_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07583__A1 _05731_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07583__B2 _01000_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08948_ _00410_ _00380_ VGND VGND VPWR VPWR _01057_ sky130_fd_sc_hd__and2_1
XANTENNA__13656__A1 _01252_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13656__B2 _01183_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08879_ _00766_ _00801_ VGND VGND VPWR VPWR _00982_ sky130_fd_sc_hd__and2b_1
X_10910_ _03201_ _03206_ VGND VGND VPWR VPWR _03207_ sky130_fd_sc_hd__xnor2_2
X_11890_ _04282_ _04102_ _04283_ VGND VGND VPWR VPWR _04284_ sky130_fd_sc_hd__nor3_1
XFILLER_0_86_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10841_ _02517_ _03130_ VGND VGND VPWR VPWR _03131_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13560_ _06071_ _06101_ VGND VGND VPWR VPWR _06103_ sky130_fd_sc_hd__nor2_1
X_10772_ _06461_ _02724_ _02727_ _02160_ VGND VGND VPWR VPWR _03055_ sky130_fd_sc_hd__a22o_1
XANTENNA__08934__A _01032_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_110 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12511_ _04958_ _04965_ _04966_ VGND VGND VPWR VPWR _04967_ sky130_fd_sc_hd__or3_1
X_13491_ _06025_ _06026_ VGND VGND VPWR VPWR _06027_ sky130_fd_sc_hd__and2_1
XFILLER_0_125_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12442_ _04886_ _04887_ _04890_ VGND VGND VPWR VPWR _04891_ sky130_fd_sc_hd__o21a_1
XFILLER_0_35_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12373_ _04813_ _04814_ VGND VGND VPWR VPWR _04815_ sky130_fd_sc_hd__xnor2_1
X_14112_ _06663_ _06665_ _06707_ VGND VGND VPWR VPWR _06708_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_50_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11324_ _03658_ _03660_ _03661_ VGND VGND VPWR VPWR _03662_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_120_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14043_ _06586_ _06633_ VGND VGND VPWR VPWR _06634_ sky130_fd_sc_hd__nor2_1
X_11255_ _03548_ _03549_ _02588_ VGND VGND VPWR VPWR _03586_ sky130_fd_sc_hd__a21o_1
X_10206_ _01995_ _02001_ _02102_ VGND VGND VPWR VPWR _02435_ sky130_fd_sc_hd__o21a_1
XANTENNA__09563__A2 _00859_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11186_ _03506_ _03509_ VGND VGND VPWR VPWR _03511_ sky130_fd_sc_hd__and2b_2
XFILLER_0_101_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12341__D _00959_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10137_ _05203_ net45 VGND VGND VPWR VPWR _02359_ sky130_fd_sc_hd__nand2_1
X_10068_ _02246_ _02247_ _01839_ VGND VGND VPWR VPWR _02283_ sky130_fd_sc_hd__and3_1
XFILLER_0_89_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13734__B _02725_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08828__B net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09005__A _06885_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13827_ _01066_ _03679_ _06396_ VGND VGND VPWR VPWR _06397_ sky130_fd_sc_hd__and3_1
XFILLER_0_58_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_767 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13758_ _06300_ _06308_ VGND VGND VPWR VPWR _06321_ sky130_fd_sc_hd__and2_1
XFILLER_0_128_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12709_ _04993_ _05031_ _04991_ VGND VGND VPWR VPWR _05185_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_127_132 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13689_ _01289_ _02730_ _06244_ VGND VGND VPWR VPWR _06245_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_128_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_664 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13583__B1 _03783_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13335__B1 _02728_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09920_ _01361_ _00159_ _02119_ _02120_ VGND VGND VPWR VPWR _02121_ sky130_fd_sc_hd__nand4_2
XFILLER_0_111_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09851_ _01633_ _01634_ _01835_ _01836_ VGND VGND VPWR VPWR _02046_ sky130_fd_sc_hd__and4_2
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08802_ _00565_ _00722_ _00727_ VGND VGND VPWR VPWR _00897_ sky130_fd_sc_hd__a21o_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09782_ _01968_ _01969_ VGND VGND VPWR VPWR _01970_ sky130_fd_sc_hd__xnor2_1
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08733_ _00817_ _00821_ VGND VGND VPWR VPWR _00822_ sky130_fd_sc_hd__xor2_1
XFILLER_0_22_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08738__B _00293_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11445__A _00262_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08664_ _00157_ _00745_ _00743_ _00583_ VGND VGND VPWR VPWR _00746_ sky130_fd_sc_hd__a31o_1
XFILLER_0_68_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__13363__C _02720_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07615_ _06032_ _06087_ VGND VGND VPWR VPWR _06098_ sky130_fd_sc_hd__xnor2_4
XTAP_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08595_ _06472_ _00257_ _00670_ _06483_ VGND VGND VPWR VPWR _00671_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_49_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07546_ _02456_ _00399_ _05335_ VGND VGND VPWR VPWR _05357_ sky130_fd_sc_hd__a21o_1
XANTENNA__08754__A _06937_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13810__A1 _02189_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13810__B2 _02188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09490__A1 _03587_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07477_ _04455_ VGND VGND VPWR VPWR _04598_ sky130_fd_sc_hd__buf_4
XFILLER_0_76_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_817 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09490__B2 _03576_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09216_ _01152_ _01349_ VGND VGND VPWR VPWR _01351_ sky130_fd_sc_hd__or2_2
XFILLER_0_63_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09147_ _01361_ _01405_ _01272_ _01211_ VGND VGND VPWR VPWR _01275_ sky130_fd_sc_hd__nand4_1
XFILLER_0_31_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09078_ _01193_ _01199_ VGND VGND VPWR VPWR _01200_ sky130_fd_sc_hd__xor2_1
XFILLER_0_32_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08029_ _07069_ _00071_ VGND VGND VPWR VPWR _00073_ sky130_fd_sc_hd__or2_1
XANTENNA__07817__B net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11040_ _03338_ _03341_ VGND VGND VPWR VPWR _03350_ sky130_fd_sc_hd__xor2_1
X_12991_ _05480_ _05483_ VGND VGND VPWR VPWR _05495_ sky130_fd_sc_hd__xor2_2
XFILLER_0_98_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11942_ _04262_ _04265_ _04339_ VGND VGND VPWR VPWR _04341_ sky130_fd_sc_hd__nor3_1
XFILLER_0_99_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12852__A2 _02306_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08367__C net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11873_ _04260_ _04262_ _04263_ _04264_ VGND VGND VPWR VPWR _04265_ sky130_fd_sc_hd__nor4_1
XFILLER_0_39_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13612_ _06157_ _06159_ VGND VGND VPWR VPWR _06160_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10824_ _01372_ _04268_ _02312_ net57 VGND VGND VPWR VPWR _03112_ sky130_fd_sc_hd__and4_1
XFILLER_0_39_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13801__A1 _02189_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13543_ _05994_ _06001_ _06053_ VGND VGND VPWR VPWR _06084_ sky130_fd_sc_hd__and3_1
XFILLER_0_39_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10755_ _00526_ _01061_ _03035_ VGND VGND VPWR VPWR _03036_ sky130_fd_sc_hd__a21o_1
XANTENNA__08284__A2 _06873_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13474_ _05992_ _06007_ VGND VGND VPWR VPWR _06008_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10686_ _05181_ _01058_ VGND VGND VPWR VPWR _02961_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10418__B _01306_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12425_ _04847_ _04870_ _04871_ VGND VGND VPWR VPWR _04872_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_113_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09495__A _00431_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12356_ _04783_ _04795_ VGND VGND VPWR VPWR _04797_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11307_ _02910_ _03633_ _03630_ VGND VGND VPWR VPWR _03644_ sky130_fd_sc_hd__nor3_1
XFILLER_0_121_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12287_ _04717_ _04720_ VGND VGND VPWR VPWR _04721_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output74_A net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14026_ _05648_ _06611_ VGND VGND VPWR VPWR _06616_ sky130_fd_sc_hd__nand2_1
X_11238_ _02978_ _02979_ VGND VGND VPWR VPWR _03568_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11169_ _03051_ _03491_ VGND VGND VPWR VPWR _03492_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10600__C _01410_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_199 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07400_ _02127_ _00322_ _03707_ _03740_ VGND VGND VPWR VPWR _03751_ sky130_fd_sc_hd__and4_1
XFILLER_0_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08380_ _00434_ _00435_ VGND VGND VPWR VPWR _00436_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07331_ _02982_ VGND VGND VPWR VPWR _02993_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_128_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07262_ _01952_ _02226_ VGND VGND VPWR VPWR _02237_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09001_ _01036_ _01039_ VGND VGND VPWR VPWR _01115_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10328__B _00373_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12246__D _01248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07193_ _01120_ _01470_ VGND VGND VPWR VPWR _01481_ sky130_fd_sc_hd__nand2_1
XFILLER_0_131_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11031__A1 net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_116 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07918__A net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11031__B2 _05027_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09903_ _02100_ _02101_ VGND VGND VPWR VPWR _02102_ sky130_fd_sc_hd__nor2_1
XANTENNA__11159__B _03480_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09834_ _02025_ _02026_ VGND VGND VPWR VPWR _02027_ sky130_fd_sc_hd__and2b_1
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10542__B1 _02728_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09765_ _01868_ _01950_ VGND VGND VPWR VPWR _01951_ sky130_fd_sc_hd__xor2_2
X_08716_ _00629_ _00802_ VGND VGND VPWR VPWR _00804_ sky130_fd_sc_hd__xnor2_1
X_09696_ _01873_ _01874_ VGND VGND VPWR VPWR _01876_ sky130_fd_sc_hd__nor2_1
XTAP_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer30 _00923_ VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__clkbuf_1
XTAP_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer41 _03378_ VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_83_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08647_ _00589_ _00592_ _00579_ VGND VGND VPWR VPWR _00728_ sky130_fd_sc_hd__o21a_1
XFILLER_0_96_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08578_ _00651_ _00652_ VGND VGND VPWR VPWR _00653_ sky130_fd_sc_hd__xnor2_1
XTAP_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07529_ _05148_ _05159_ VGND VGND VPWR VPWR _05170_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08266__A2 _00310_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10540_ _00294_ _02169_ VGND VGND VPWR VPWR _02800_ sky130_fd_sc_hd__nand2_1
XFILLER_0_106_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09215__A1 _01155_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10471_ _02723_ VGND VGND VPWR VPWR _02724_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12210_ _04633_ _04635_ VGND VGND VPWR VPWR _04636_ sky130_fd_sc_hd__or2_1
X_13190_ _05705_ _05706_ VGND VGND VPWR VPWR _05714_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08650__C net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12141_ _04475_ _04476_ VGND VGND VPWR VPWR _04560_ sky130_fd_sc_hd__nor2_1
XFILLER_0_102_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12072_ _04473_ _04483_ VGND VGND VPWR VPWR _04484_ sky130_fd_sc_hd__nor2_1
X_11023_ _03326_ _03328_ _03330_ VGND VGND VPWR VPWR _03331_ sky130_fd_sc_hd__o21a_1
XANTENNA__08659__A _03938_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10701__B _01059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12974_ _05475_ VGND VGND VPWR VPWR _05476_ sky130_fd_sc_hd__inv_2
X_11925_ _04287_ _04321_ VGND VGND VPWR VPWR _04322_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_87_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output112_A net112 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07701__A1 net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07701__B2 net1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_840 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11856_ _04245_ _02692_ _02689_ VGND VGND VPWR VPWR _04247_ sky130_fd_sc_hd__a21o_1
XFILLER_0_129_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12589__A1 _00745_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10807_ _03089_ VGND VGND VPWR VPWR _03094_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11787_ _04164_ _04170_ VGND VGND VPWR VPWR _04171_ sky130_fd_sc_hd__xor2_1
XFILLER_0_82_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13526_ _06040_ _06064_ VGND VGND VPWR VPWR _06066_ sky130_fd_sc_hd__xor2_1
XANTENNA__08544__D _00613_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10738_ _03015_ _02758_ _02720_ _00399_ VGND VGND VPWR VPWR _03018_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13457_ _05983_ _05987_ VGND VGND VPWR VPWR _05990_ sky130_fd_sc_hd__or2_1
X_10669_ _05181_ _01411_ _02940_ _02941_ VGND VGND VPWR VPWR _02942_ sky130_fd_sc_hd__a31o_1
XFILLER_0_88_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12408_ _04059_ _01272_ _04852_ _04853_ VGND VGND VPWR VPWR _04854_ sky130_fd_sc_hd__a31o_1
XFILLER_0_106_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13388_ _05384_ _05391_ VGND VGND VPWR VPWR _05915_ sky130_fd_sc_hd__and2_1
Xoutput106 net106 VGND VGND VPWR VPWR prod[47] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput117 net117 VGND VGND VPWR VPWR prod[57] sky130_fd_sc_hd__clkbuf_4
Xoutput128 net128 VGND VGND VPWR VPWR prod[9] sky130_fd_sc_hd__buf_2
X_12339_ _00755_ _01260_ _01507_ _01369_ VGND VGND VPWR VPWR _04778_ sky130_fd_sc_hd__nand4_2
XFILLER_0_121_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10772__B1 _02727_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14009_ _06521_ _06532_ VGND VGND VPWR VPWR _06597_ sky130_fd_sc_hd__and2b_1
XANTENNA__13475__A _02856_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07880_ _00891_ net37 _06953_ _06952_ VGND VGND VPWR VPWR _07009_ sky130_fd_sc_hd__a31o_1
XFILLER_0_128_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13194__B _05704_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09550_ _01713_ _01715_ VGND VGND VPWR VPWR _01716_ sky130_fd_sc_hd__xor2_2
XANTENNA__08719__D _04873_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08501_ _00350_ _00568_ _00372_ _00411_ VGND VGND VPWR VPWR _00569_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_77_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09481_ _01636_ _01640_ VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__xor2_4
XFILLER_0_144_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09693__A1 _05192_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08432_ _00469_ _00492_ VGND VGND VPWR VPWR _00493_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_144_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08363_ _00333_ _00416_ VGND VGND VPWR VPWR _00417_ sky130_fd_sc_hd__nand2_2
XFILLER_0_19_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_759 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07314_ _02631_ _02795_ VGND VGND VPWR VPWR _02806_ sky130_fd_sc_hd__nor2_1
X_08294_ _00340_ _00341_ VGND VGND VPWR VPWR _00342_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07245_ _00989_ VGND VGND VPWR VPWR _02051_ sky130_fd_sc_hd__buf_4
XFILLER_0_73_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08751__B _00703_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11004__A1 _04598_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07648__A _05588_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11004__B2 _05203_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07176_ _01197_ VGND VGND VPWR VPWR _01295_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11555__A2 _01564_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_845 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08479__A _00399_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09817_ _00530_ _02008_ VGND VGND VPWR VPWR _02009_ sky130_fd_sc_hd__nand2_1
X_09748_ net53 VGND VGND VPWR VPWR _01933_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__09133__B1 _03938_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09679_ _01855_ _01856_ VGND VGND VPWR VPWR _01857_ sky130_fd_sc_hd__nor2_1
XTAP_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12729__A _05193_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08926__B _00871_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11710_ _00258_ _00915_ VGND VGND VPWR VPWR _04086_ sky130_fd_sc_hd__nand2_1
XTAP_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_158 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12690_ _04910_ _05163_ VGND VGND VPWR VPWR _05164_ sky130_fd_sc_hd__and2_1
XTAP_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11641_ _03735_ _03843_ VGND VGND VPWR VPWR _04010_ sky130_fd_sc_hd__or2_1
XANTENNA__11352__B _03680_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_342 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11572_ _03924_ _03932_ _03933_ VGND VGND VPWR VPWR _03934_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_80_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13311_ _05786_ _05802_ _05831_ _05832_ VGND VGND VPWR VPWR _05833_ sky130_fd_sc_hd__a31o_2
XFILLER_0_18_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput19 a[26] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__buf_4
X_10523_ _02754_ _02780_ VGND VGND VPWR VPWR _02781_ sky130_fd_sc_hd__or2_1
XFILLER_0_64_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08661__B _00742_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_135_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13242_ _05572_ _05568_ _05570_ VGND VGND VPWR VPWR _05767_ sky130_fd_sc_hd__nand3_1
XANTENNA__07558__A _05478_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10454_ _02482_ VGND VGND VPWR VPWR _02706_ sky130_fd_sc_hd__inv_2
XANTENNA__11546__A2 _02120_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12743__A1 _01953_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13173_ _05683_ _05689_ VGND VGND VPWR VPWR _05695_ sky130_fd_sc_hd__xor2_2
XANTENNA__08411__A2 _07004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10385_ _02418_ _02629_ VGND VGND VPWR VPWR _02630_ sky130_fd_sc_hd__nor2_1
XFILLER_0_103_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12124_ _04525_ _04527_ VGND VGND VPWR VPWR _04541_ sky130_fd_sc_hd__nor2_1
XANTENNA__09773__A net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12055_ _04461_ _04464_ VGND VGND VPWR VPWR _04465_ sky130_fd_sc_hd__nand2_2
XANTENNA__10506__B1 _02726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11006_ _03308_ _03311_ VGND VGND VPWR VPWR _03313_ sky130_fd_sc_hd__nor2_1
XANTENNA__13445__D _02722_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08539__D _00608_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13742__B _02858_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12957_ _04534_ _04535_ VGND VGND VPWR VPWR _05458_ sky130_fd_sc_hd__or2_1
XFILLER_0_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11543__A _03521_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11908_ _04291_ _04302_ VGND VGND VPWR VPWR _04304_ sky130_fd_sc_hd__or2_1
XTAP_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12888_ _00379_ _03678_ _05226_ VGND VGND VPWR VPWR _05382_ sky130_fd_sc_hd__and3_1
XFILLER_0_75_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11839_ _03070_ _01955_ _03686_ _02456_ VGND VGND VPWR VPWR _04228_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_74_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10037__A2 _01473_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_720 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13509_ _06031_ _06046_ VGND VGND VPWR VPWR _06047_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_55_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09667__B _00859_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12374__A _00389_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08571__B _06966_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11537__A2 _01178_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07187__B _01405_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08981_ _01086_ _01092_ VGND VGND VPWR VPWR _01093_ sky130_fd_sc_hd__xor2_1
X_07932_ _07059_ _07060_ net44 net7 VGND VGND VPWR VPWR _07061_ sky130_fd_sc_hd__and4bb_1
XANTENNA__11718__A _00263_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11437__B _03785_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07863_ _06384_ _06990_ _06615_ VGND VGND VPWR VPWR _06992_ sky130_fd_sc_hd__o21ai_1
X_09602_ _01771_ _01772_ VGND VGND VPWR VPWR _01773_ sky130_fd_sc_hd__or2_2
X_07794_ _06921_ _06922_ VGND VGND VPWR VPWR _06923_ sky130_fd_sc_hd__nor2_1
X_09533_ _01663_ _01696_ VGND VGND VPWR VPWR _01697_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07931__A net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09464_ _01614_ _01621_ VGND VGND VPWR VPWR _01622_ sky130_fd_sc_hd__xor2_2
XFILLER_0_38_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08415_ _00471_ _00473_ VGND VGND VPWR VPWR _00474_ sky130_fd_sc_hd__and2_1
XFILLER_0_65_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09395_ _01545_ VGND VGND VPWR VPWR _01546_ sky130_fd_sc_hd__buf_2
XFILLER_0_46_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08346_ _00387_ _00396_ _00398_ VGND VGND VPWR VPWR _00400_ sky130_fd_sc_hd__or3_1
XFILLER_0_34_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08277_ _00321_ _00323_ VGND VGND VPWR VPWR _00324_ sky130_fd_sc_hd__nor2_2
XFILLER_0_62_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07228_ _01219_ _01438_ _01842_ _01186_ VGND VGND VPWR VPWR _01864_ sky130_fd_sc_hd__o31ai_1
XANTENNA__07378__A _03499_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07809__C _06937_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07159_ _00880_ net59 _00945_ _00934_ VGND VGND VPWR VPWR _01109_ sky130_fd_sc_hd__a31o_1
XFILLER_0_30_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10170_ _02393_ _02394_ VGND VGND VPWR VPWR _02395_ sky130_fd_sc_hd__and2_1
XANTENNA__13827__B _03679_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13860_ _06416_ _06431_ _06432_ VGND VGND VPWR VPWR _06433_ sky130_fd_sc_hd__and3_1
XFILLER_0_88_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12811_ _05108_ _05114_ _05296_ VGND VGND VPWR VPWR _05297_ sky130_fd_sc_hd__a21o_1
X_13791_ _06292_ _06312_ VGND VGND VPWR VPWR _06357_ sky130_fd_sc_hd__nor2_1
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12742_ _00779_ _01953_ _02134_ _00784_ VGND VGND VPWR VPWR _05221_ sky130_fd_sc_hd__a22o_1
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12178__B _04600_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12673_ _05141_ _05142_ _05144_ VGND VGND VPWR VPWR _05145_ sky130_fd_sc_hd__nor3_1
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11624_ _03980_ _03977_ VGND VGND VPWR VPWR _03991_ sky130_fd_sc_hd__nand2_1
XTAP_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09768__A _01954_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08672__A _03894_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11555_ _00486_ _01564_ _03913_ _03914_ _01247_ VGND VGND VPWR VPWR _03915_ sky130_fd_sc_hd__a32o_1
XANTENNA__11810__B _03750_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08391__B _04026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10506_ _00636_ _02721_ _02726_ _00526_ VGND VGND VPWR VPWR _02763_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08822__D net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11486_ _03789_ _03790_ _03800_ _03838_ VGND VGND VPWR VPWR _03840_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_12_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13225_ _05680_ _05743_ _05751_ VGND VGND VPWR VPWR _05752_ sky130_fd_sc_hd__o21ba_1
X_10437_ _02683_ _02687_ VGND VGND VPWR VPWR _02688_ sky130_fd_sc_hd__and2b_1
XFILLER_0_110_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13156_ _05668_ _05671_ _05675_ VGND VGND VPWR VPWR _05677_ sky130_fd_sc_hd__o21a_1
XFILLER_0_103_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10368_ _02407_ _02611_ VGND VGND VPWR VPWR _02612_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_798 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12641__B _02857_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12107_ _04503_ _04514_ VGND VGND VPWR VPWR _04523_ sky130_fd_sc_hd__and2_2
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13087_ _05453_ _05471_ VGND VGND VPWR VPWR _05601_ sky130_fd_sc_hd__nor2_1
X_10299_ _02534_ _02535_ VGND VGND VPWR VPWR _02536_ sky130_fd_sc_hd__nand2_1
X_12038_ _04445_ _04446_ VGND VGND VPWR VPWR _04447_ sky130_fd_sc_hd__xnor2_2
XANTENNA__07454__C _00366_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13692__A2 _02736_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13989_ _06556_ _06559_ VGND VGND VPWR VPWR _06575_ sky130_fd_sc_hd__and2b_1
XFILLER_0_34_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08320__A1 _00352_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_854 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08200_ _00202_ _00243_ VGND VGND VPWR VPWR _00244_ sky130_fd_sc_hd__nor2_4
XFILLER_0_8_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09180_ _01027_ _01030_ _01159_ VGND VGND VPWR VPWR _01311_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_56_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08582__A _00543_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08131_ _00172_ _00174_ VGND VGND VPWR VPWR _00175_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_56_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08062_ _06472_ _06885_ _00103_ _00104_ VGND VGND VPWR VPWR _00106_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_43_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08387__A1 _04081_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11448__A _00263_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08964_ _01076_ net47 _00959_ _03587_ VGND VGND VPWR VPWR _01074_ sky130_fd_sc_hd__a22o_1
X_07915_ _06916_ _06919_ _07043_ VGND VGND VPWR VPWR _07044_ sky130_fd_sc_hd__a21o_1
X_08895_ _00508_ _00158_ _00807_ _00809_ VGND VGND VPWR VPWR _00999_ sky130_fd_sc_hd__a211o_1
X_07846_ _06872_ _06880_ _06974_ VGND VGND VPWR VPWR _06975_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10497__A2 _02721_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07777_ net33 net7 VGND VGND VPWR VPWR _06906_ sky130_fd_sc_hd__and2_1
XANTENNA__09639__A1 _00300_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09516_ _01535_ _01676_ VGND VGND VPWR VPWR _01679_ sky130_fd_sc_hd__or2_1
XANTENNA__11446__A1 _00262_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11446__B2 _00263_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07811__D net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09447_ _01599_ _01603_ VGND VGND VPWR VPWR _01604_ sky130_fd_sc_hd__xnor2_1
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11911__A _06626_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09378_ _01501_ _01526_ VGND VGND VPWR VPWR _01528_ sky130_fd_sc_hd__and2_1
XFILLER_0_35_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08329_ _00380_ VGND VGND VPWR VPWR _00381_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_46_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11340_ _03678_ VGND VGND VPWR VPWR _03679_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_15_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11271_ _03595_ _03603_ VGND VGND VPWR VPWR _03604_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13010_ _05512_ _05513_ _05514_ _05515_ VGND VGND VPWR VPWR _05516_ sky130_fd_sc_hd__and4_1
X_10222_ _02450_ _01564_ _02029_ _02448_ VGND VGND VPWR VPWR _02452_ sky130_fd_sc_hd__and4b_1
XANTENNA__07836__A _06964_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10185__A1 _06821_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10185__B2 _03499_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11358__A _03680_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10153_ _02349_ _02375_ VGND VGND VPWR VPWR _02376_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_100_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10084_ _02167_ _02174_ VGND VGND VPWR VPWR _02300_ sky130_fd_sc_hd__or2b_1
X_13912_ _06235_ _06489_ VGND VGND VPWR VPWR _06490_ sky130_fd_sc_hd__and2_1
X_13843_ _06386_ _06411_ _06413_ VGND VGND VPWR VPWR _06414_ sky130_fd_sc_hd__o21a_1
XFILLER_0_97_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10986_ _03286_ VGND VGND VPWR VPWR _03291_ sky130_fd_sc_hd__inv_2
X_13774_ _06332_ _06333_ _06337_ VGND VGND VPWR VPWR _06338_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_84_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12339__D _01369_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12725_ _05198_ _05201_ VGND VGND VPWR VPWR _05202_ sky130_fd_sc_hd__and2_1
XFILLER_0_128_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12656_ _05089_ _05085_ VGND VGND VPWR VPWR _05127_ sky130_fd_sc_hd__or2_1
XFILLER_0_127_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11607_ _03966_ _03972_ VGND VGND VPWR VPWR _03973_ sky130_fd_sc_hd__xnor2_2
XANTENNA__11540__B _06874_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12587_ _00915_ _01412_ _05048_ _05050_ VGND VGND VPWR VPWR _05051_ sky130_fd_sc_hd__a31o_1
XFILLER_0_52_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11538_ _03895_ _03896_ _03510_ _01564_ VGND VGND VPWR VPWR _03897_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_111_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_cap138 _03504_ VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__buf_1
X_11469_ _03816_ _03820_ VGND VGND VPWR VPWR _03821_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12652__A _00390_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08369__B2 _01306_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07746__A _06874_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13208_ _05715_ _05724_ VGND VGND VPWR VPWR _05734_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14188_ _06613_ _06617_ VGND VGND VPWR VPWR _06787_ sky130_fd_sc_hd__nor2_2
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13139_ _05212_ _05657_ VGND VGND VPWR VPWR _05658_ sky130_fd_sc_hd__nor2_1
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07700_ _06827_ _06828_ VGND VGND VPWR VPWR _06829_ sky130_fd_sc_hd__nor2_1
XANTENNA__13483__A _02858_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08680_ _00729_ _00763_ VGND VGND VPWR VPWR _00764_ sky130_fd_sc_hd__xnor2_4
XANTENNA__07344__A2 net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07631_ _06186_ _06252_ VGND VGND VPWR VPWR _06274_ sky130_fd_sc_hd__nor2_1
XANTENNA__07481__A _00300_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07562_ _05434_ _05500_ _03169_ VGND VGND VPWR VPWR _05533_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_88_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12625__B1 _02306_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09301_ _00557_ _01167_ _01441_ _01442_ VGND VGND VPWR VPWR _01443_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_146_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07493_ _03037_ _04763_ VGND VGND VPWR VPWR _04774_ sky130_fd_sc_hd__and2_1
XFILLER_0_61_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09232_ net47 VGND VGND VPWR VPWR _01368_ sky130_fd_sc_hd__buf_2
XFILLER_0_145_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09201__A _06965_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09163_ _01291_ VGND VGND VPWR VPWR _01292_ sky130_fd_sc_hd__inv_2
XANTENNA__12209__A1_N _00379_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13050__B1 _05559_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08114_ net7 VGND VGND VPWR VPWR _00158_ sky130_fd_sc_hd__clkbuf_4
X_09094_ _00910_ _01216_ VGND VGND VPWR VPWR _01217_ sky130_fd_sc_hd__nand2_1
XANTENNA__07359__C _02664_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10066__B _01867_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08045_ _00086_ _00087_ _00088_ VGND VGND VPWR VPWR _00089_ sky130_fd_sc_hd__or3_4
XFILLER_0_102_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11903__A2 _03678_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09996_ _01904_ _02202_ VGND VGND VPWR VPWR _02205_ sky130_fd_sc_hd__nand2_1
XANTENNA__07583__A2 _00628_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08947_ _01050_ _01052_ VGND VGND VPWR VPWR _01056_ sky130_fd_sc_hd__and2_4
XANTENNA__13656__A2 _02766_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_816 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08878_ _00976_ _00980_ VGND VGND VPWR VPWR _00981_ sky130_fd_sc_hd__xnor2_2
X_07829_ _01120_ _06744_ VGND VGND VPWR VPWR _06958_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10840_ _03127_ _03128_ VGND VGND VPWR VPWR _03130_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_39_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10771_ _02160_ _06461_ _02724_ _02727_ VGND VGND VPWR VPWR _03054_ sky130_fd_sc_hd__and4_1
XFILLER_0_67_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12510_ _04947_ _04951_ VGND VGND VPWR VPWR _04966_ sky130_fd_sc_hd__xor2_1
XFILLER_0_136_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13490_ _01062_ _03699_ _06011_ _06013_ VGND VGND VPWR VPWR _06026_ sky130_fd_sc_hd__a211o_1
XFILLER_0_94_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12441_ _04886_ _04887_ _04889_ VGND VGND VPWR VPWR _04890_ sky130_fd_sc_hd__a21o_1
XFILLER_0_136_166 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08048__B1 _06875_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_805 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12372_ _00914_ _00457_ VGND VGND VPWR VPWR _04814_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14111_ _06705_ _06706_ VGND VGND VPWR VPWR _06707_ sky130_fd_sc_hd__xnor2_1
X_11323_ _02917_ _03657_ _03655_ VGND VGND VPWR VPWR _03661_ sky130_fd_sc_hd__or3_1
XFILLER_0_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_860 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09548__B1 _01500_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07566__A _02664_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11254_ _03551_ _03552_ _03584_ VGND VGND VPWR VPWR _03585_ sky130_fd_sc_hd__a21o_1
XFILLER_0_120_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14042_ _06629_ _06577_ net135 VGND VGND VPWR VPWR _06633_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_120_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10205_ _02431_ _02432_ VGND VGND VPWR VPWR _02433_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11185_ net138 _03505_ _03508_ VGND VGND VPWR VPWR _03509_ sky130_fd_sc_hd__a21o_1
XFILLER_0_66_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10136_ _01506_ _02224_ _02356_ VGND VGND VPWR VPWR _02358_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_100_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09781__A _01744_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10067_ _02268_ _02281_ VGND VGND VPWR VPWR _02282_ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10330__A1 _05027_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09005__B _00294_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13826_ _00460_ _03683_ _06388_ _06387_ _01955_ VGND VGND VPWR VPWR _06396_ sky130_fd_sc_hd__a32o_1
XFILLER_0_57_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_735 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13757_ _06316_ _06319_ VGND VGND VPWR VPWR _06320_ sky130_fd_sc_hd__nand2_1
X_10969_ _03271_ VGND VGND VPWR VPWR _03272_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_779 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12708_ _04991_ _04993_ _05031_ VGND VGND VPWR VPWR _05184_ sky130_fd_sc_hd__and3_1
XFILLER_0_45_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13688_ _02090_ _02725_ VGND VGND VPWR VPWR _06244_ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09021__A _06964_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12639_ _05106_ _05107_ VGND VGND VPWR VPWR _05108_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_199 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13583__A1 _03785_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_142_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13583__B2 _02856_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_158 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13335__A1 _00745_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13335__B2 _00914_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09850_ _01833_ _02044_ VGND VGND VPWR VPWR _02045_ sky130_fd_sc_hd__xor2_4
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08801_ _00894_ _00896_ VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__xor2_2
XANTENNA__09691__A _05181_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09781_ _01744_ net20 VGND VGND VPWR VPWR _01969_ sky130_fd_sc_hd__nand2_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08732_ _00262_ _00818_ _00820_ VGND VGND VPWR VPWR _00821_ sky130_fd_sc_hd__and3_1
XANTENNA__10630__A _00818_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09711__B1 _01505_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08663_ _00741_ VGND VGND VPWR VPWR _00745_ sky130_fd_sc_hd__buf_4
XANTENNA__11445__B _00263_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08100__A _00143_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07614_ _05999_ _06010_ VGND VGND VPWR VPWR _06087_ sky130_fd_sc_hd__xor2_2
XFILLER_0_95_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08594_ _00258_ VGND VGND VPWR VPWR _00670_ sky130_fd_sc_hd__buf_4
XTAP_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07545_ _02335_ _00399_ _05335_ VGND VGND VPWR VPWR _05346_ sky130_fd_sc_hd__and3_1
XFILLER_0_49_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08754__B _00844_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13810__A2 _01955_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11461__A _03532_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07476_ _04565_ _04576_ VGND VGND VPWR VPWR _04587_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09215_ _01155_ _01156_ _01154_ VGND VGND VPWR VPWR _01349_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11180__B _03501_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09146_ _01295_ _01272_ _01211_ _01405_ VGND VGND VPWR VPWR _01274_ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09077_ _01196_ _01198_ VGND VGND VPWR VPWR _01199_ sky130_fd_sc_hd__nor2_1
XFILLER_0_114_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07386__A _03576_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08028_ _07069_ _00071_ VGND VGND VPWR VPWR _00072_ sky130_fd_sc_hd__nand2_1
X_09979_ _06637_ _01400_ _01892_ _01893_ VGND VGND VPWR VPWR _02186_ sky130_fd_sc_hd__a31o_1
XANTENNA__10540__A _00294_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12990_ _04581_ _05442_ VGND VGND VPWR VPWR _05494_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_99_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11941_ _04262_ net146 _04339_ VGND VGND VPWR VPWR _04340_ sky130_fd_sc_hd__o21a_1
XANTENNA__10312__A1 _01369_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08367__D net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11872_ _07004_ _01780_ _04261_ VGND VGND VPWR VPWR _04264_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11357__A1_N _01312_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13611_ _06150_ _06158_ VGND VGND VPWR VPWR _06159_ sky130_fd_sc_hd__nor2_1
X_10823_ _01339_ net54 _03109_ _03110_ VGND VGND VPWR VPWR _03111_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_39_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13801__A2 _03686_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_420 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13542_ _06048_ _06073_ _06082_ VGND VGND VPWR VPWR _06083_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_27_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10754_ _00399_ _02759_ _03033_ VGND VGND VPWR VPWR _03035_ sky130_fd_sc_hd__and3_1
XFILLER_0_48_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13473_ _06005_ _06006_ VGND VGND VPWR VPWR _06007_ sky130_fd_sc_hd__nor2_1
X_10685_ _02956_ _02958_ VGND VGND VPWR VPWR _02959_ sky130_fd_sc_hd__and2_1
XFILLER_0_124_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10418__C net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12424_ _04841_ _04844_ _04846_ VGND VGND VPWR VPWR _04871_ sky130_fd_sc_hd__and3_1
XFILLER_0_23_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10379__A1 _00475_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09495__B _04169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12355_ _04778_ _04782_ _04781_ VGND VGND VPWR VPWR _04795_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_121_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11306_ _03637_ _03641_ VGND VGND VPWR VPWR _03643_ sky130_fd_sc_hd__or2_1
X_12286_ _00380_ _01956_ _04718_ VGND VGND VPWR VPWR _04720_ sky130_fd_sc_hd__a21o_1
XFILLER_0_121_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11237_ _03563_ _03566_ VGND VGND VPWR VPWR _03567_ sky130_fd_sc_hd__and2b_1
XANTENNA__12352__D _01369_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14025_ _05810_ _05811_ _05812_ _05835_ VGND VGND VPWR VPWR _06614_ sky130_fd_sc_hd__a31o_1
XFILLER_0_120_397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_output67_A net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11168_ _03003_ _03050_ VGND VGND VPWR VPWR _03491_ sky130_fd_sc_hd__and2_1
XFILLER_0_93_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10119_ _02195_ _02338_ VGND VGND VPWR VPWR _02339_ sky130_fd_sc_hd__xor2_1
X_11099_ _00635_ _01066_ _03414_ _07040_ VGND VGND VPWR VPWR _03415_ sky130_fd_sc_hd__a22oi_1
XANTENNA__13464__C _02735_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10600__D _02158_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13809_ _02187_ _02189_ _01954_ _03686_ VGND VGND VPWR VPWR _06377_ sky130_fd_sc_hd__and4_1
XFILLER_0_133_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07330_ _02971_ VGND VGND VPWR VPWR _02982_ sky130_fd_sc_hd__buf_4
XFILLER_0_18_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07261_ _01908_ _01919_ VGND VGND VPWR VPWR _02226_ sky130_fd_sc_hd__xor2_1
XFILLER_0_6_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09000_ _01034_ _01040_ _01032_ VGND VGND VPWR VPWR _01114_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_26_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07192_ _00661_ VGND VGND VPWR VPWR _01470_ sky130_fd_sc_hd__buf_4
XFILLER_0_14_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11031__A2 _00782_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07918__B net61 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09902_ _02098_ _02099_ VGND VGND VPWR VPWR _02101_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09833_ _07004_ _00390_ _02024_ VGND VGND VPWR VPWR _02026_ sky130_fd_sc_hd__a21o_1
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10542__A1 _03004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10542__B2 _00388_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09764_ _01947_ _01948_ _01949_ VGND VGND VPWR VPWR _01950_ sky130_fd_sc_hd__nor3_2
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10360__A _06733_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08715_ _00766_ _00801_ VGND VGND VPWR VPWR _00802_ sky130_fd_sc_hd__xnor2_1
X_09695_ _02960_ _04367_ _04180_ _04191_ VGND VGND VPWR VPWR _01874_ sky130_fd_sc_hd__and4_1
Xrebuffer20 _06934_ VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__buf_1
XTAP_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer31 _00923_ VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__clkbuf_2
XTAP_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08646_ _00718_ _00719_ VGND VGND VPWR VPWR _00727_ sky130_fd_sc_hd__and2_2
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07171__B1 _01208_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08577_ _00340_ _00539_ _00538_ VGND VGND VPWR VPWR _00652_ sky130_fd_sc_hd__o21ba_1
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07528_ _05115_ _05137_ _04345_ VGND VGND VPWR VPWR _05159_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_76_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07459_ net58 net163 net31 net32 VGND VGND VPWR VPWR _04400_ sky130_fd_sc_hd__and4_1
XFILLER_0_119_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10470_ _02312_ VGND VGND VPWR VPWR _02723_ sky130_fd_sc_hd__buf_2
XFILLER_0_91_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09215__A2 _01156_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09129_ _02138_ _00322_ _01179_ _01254_ VGND VGND VPWR VPWR _01255_ sky130_fd_sc_hd__nand4_4
XFILLER_0_115_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12140_ _02596_ _02644_ _02693_ VGND VGND VPWR VPWR _04559_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_114_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08650__D _00730_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08005__A _01044_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12071_ _04479_ _04481_ _04482_ VGND VGND VPWR VPWR _04483_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11022_ _03321_ _03329_ VGND VGND VPWR VPWR _03330_ sky130_fd_sc_hd__nor2_1
XANTENNA__12286__A1 _00380_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12973_ _05433_ _05447_ VGND VGND VPWR VPWR _05475_ sky130_fd_sc_hd__xor2_2
X_11924_ _04289_ _04320_ VGND VGND VPWR VPWR _04321_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_86_115 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07701__A2 net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_852 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11855_ _02683_ _02687_ VGND VGND VPWR VPWR _04245_ sky130_fd_sc_hd__or2b_1
XFILLER_0_86_159 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_output105_A net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12589__A2 _01412_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10806_ _03082_ _03091_ VGND VGND VPWR VPWR _03093_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11786_ _02454_ _02659_ _04167_ _04168_ VGND VGND VPWR VPWR _04170_ sky130_fd_sc_hd__o31a_1
XFILLER_0_82_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12994__C1 _02008_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13525_ _06062_ _06063_ VGND VGND VPWR VPWR _06064_ sky130_fd_sc_hd__nor2_1
X_10737_ _00399_ _03015_ _02758_ _02721_ VGND VGND VPWR VPWR _03017_ sky130_fd_sc_hd__nand4_1
XFILLER_0_82_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13456_ _05983_ _05987_ VGND VGND VPWR VPWR _05989_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_387 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_410 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10668_ _02982_ _05192_ _01546_ _02156_ VGND VGND VPWR VPWR _02941_ sky130_fd_sc_hd__and4_1
XFILLER_0_70_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12407_ _00373_ _00782_ _00413_ _00571_ VGND VGND VPWR VPWR _04853_ sky130_fd_sc_hd__and4_1
XFILLER_0_112_117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13387_ _05383_ _05392_ VGND VGND VPWR VPWR _05914_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10599_ _02853_ _02864_ VGND VGND VPWR VPWR _02865_ sky130_fd_sc_hd__xor2_1
XFILLER_0_51_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput107 net107 VGND VGND VPWR VPWR prod[48] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_112_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput118 net118 VGND VGND VPWR VPWR prod[58] sky130_fd_sc_hd__clkbuf_4
X_12338_ _04772_ _04776_ VGND VGND VPWR VPWR _04777_ sky130_fd_sc_hd__nor2_1
XFILLER_0_50_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10772__A1 _06461_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12269_ _04638_ _04700_ VGND VGND VPWR VPWR _04701_ sky130_fd_sc_hd__xnor2_1
X_14008_ net132 _06587_ _06592_ _06595_ VGND VGND VPWR VPWR _06596_ sky130_fd_sc_hd__o31a_2
XFILLER_0_128_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08500_ _00371_ VGND VGND VPWR VPWR _00568_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09480_ _01637_ net131 _01433_ _01639_ VGND VGND VPWR VPWR _01640_ sky130_fd_sc_hd__a31o_2
XANTENNA__09693__A2 _00373_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08431_ _00490_ _00491_ VGND VGND VPWR VPWR _00492_ sky130_fd_sc_hd__nor2_2
XFILLER_0_59_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08362_ _00415_ VGND VGND VPWR VPWR _00416_ sky130_fd_sc_hd__buf_4
XFILLER_0_58_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07313_ net153 _02784_ VGND VGND VPWR VPWR _02795_ sky130_fd_sc_hd__xnor2_1
X_08293_ _00098_ _00339_ VGND VGND VPWR VPWR _00341_ sky130_fd_sc_hd__or2_1
XANTENNA__12835__A _00916_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07244_ _02029_ VGND VGND VPWR VPWR _02040_ sky130_fd_sc_hd__buf_4
XFILLER_0_33_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_242 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07175_ _01076_ VGND VGND VPWR VPWR _01284_ sky130_fd_sc_hd__buf_4
XFILLER_0_131_426 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__07664__A _06494_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13701__A1 _02426_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__08479__B _00544_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09816_ _01188_ VGND VGND VPWR VPWR _02008_ sky130_fd_sc_hd__buf_4
XANTENNA__10090__A _01383_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09747_ _01661_ _01931_ VGND VGND VPWR VPWR _01932_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09133__A1 _05456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09133__B2 _05467_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08495__A _00439_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07144__B1 net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09678_ _01838_ _01854_ VGND VGND VPWR VPWR _01856_ sky130_fd_sc_hd__nor2_1
XFILLER_0_69_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08629_ _00466_ _00524_ _00708_ VGND VGND VPWR VPWR _00709_ sky130_fd_sc_hd__o21a_1
XTAP_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11640_ _03862_ _04008_ VGND VGND VPWR VPWR _04009_ sky130_fd_sc_hd__and2b_1
XTAP_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11571_ _03917_ _03922_ _03923_ VGND VGND VPWR VPWR _03933_ sky130_fd_sc_hd__o21a_1
XFILLER_0_64_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13310_ _05805_ _05831_ VGND VGND VPWR VPWR _05832_ sky130_fd_sc_hd__and2_1
XFILLER_0_52_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10522_ _02753_ _02749_ VGND VGND VPWR VPWR _02780_ sky130_fd_sc_hd__and2b_1
XFILLER_0_107_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10453_ _02592_ _02593_ _02703_ VGND VGND VPWR VPWR _02705_ sky130_fd_sc_hd__a21o_1
X_13241_ _05562_ _05766_ VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__xnor2_4
XANTENNA__07558__B _01383_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09076__A1_N _01996_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10384_ _02627_ _02628_ VGND VGND VPWR VPWR _02629_ sky130_fd_sc_hd__nand2_1
X_13172_ _05682_ _05693_ VGND VGND VPWR VPWR _05694_ sky130_fd_sc_hd__xor2_4
XFILLER_0_103_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12123_ _04539_ VGND VGND VPWR VPWR _04540_ sky130_fd_sc_hd__inv_2
XANTENNA__13576__A _02855_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12054_ _04462_ _04463_ VGND VGND VPWR VPWR _04464_ sky130_fd_sc_hd__nor2_1
XANTENNA__10506__A1 _00636_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10506__B2 _00526_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11005_ _03309_ _03310_ VGND VGND VPWR VPWR _03311_ sky130_fd_sc_hd__or2_1
XFILLER_0_74_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__07383__B1 _00519_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12956_ _05426_ _05429_ VGND VGND VPWR VPWR _05457_ sky130_fd_sc_hd__nor2_1
X_11907_ _04291_ _04302_ VGND VGND VPWR VPWR _04303_ sky130_fd_sc_hd__nand2_1
XANTENNA__11543__B _01960_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12887_ _05226_ _05227_ VGND VGND VPWR VPWR _05381_ sky130_fd_sc_hd__or2b_1
XFILLER_0_23_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11838_ _04223_ _04226_ VGND VGND VPWR VPWR _04227_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_855 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11769_ _02007_ _01564_ _02649_ _02648_ _01178_ VGND VGND VPWR VPWR _04151_ sky130_fd_sc_hd__a32o_1
XFILLER_0_126_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_743 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13508_ _06044_ _06045_ VGND VGND VPWR VPWR _06046_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12374__B _00392_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08571__C _00095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_140_201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13439_ _01181_ _01250_ _02721_ _02726_ VGND VGND VPWR VPWR _05970_ sky130_fd_sc_hd__and4_1
XFILLER_0_140_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09964__A _02168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08980_ _01090_ _01091_ VGND VGND VPWR VPWR _01092_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07931_ net58 _00716_ net6 net5 VGND VGND VPWR VPWR _07060_ sky130_fd_sc_hd__and4_1
XANTENNA__11718__B _01600_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07862_ _06384_ _06615_ _06990_ VGND VGND VPWR VPWR _06991_ sky130_fd_sc_hd__or3_1
X_09601_ _01302_ _01620_ _01770_ VGND VGND VPWR VPWR _01772_ sky130_fd_sc_hd__o21a_1
X_07793_ _05148_ _06920_ VGND VGND VPWR VPWR _06922_ sky130_fd_sc_hd__and2_1
X_09532_ _01692_ _01695_ VGND VGND VPWR VPWR _01696_ sky130_fd_sc_hd__xnor2_2
X_09463_ _01302_ _01620_ VGND VGND VPWR VPWR _01621_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_66_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08414_ _00472_ VGND VGND VPWR VPWR _00473_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09394_ net51 VGND VGND VPWR VPWR _01545_ sky130_fd_sc_hd__buf_2
XFILLER_0_93_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08345_ _00352_ _00397_ VGND VGND VPWR VPWR _00398_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_74_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11630__C1 _01958_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08276_ _00319_ _00320_ VGND VGND VPWR VPWR _00323_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_724 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07227_ _01186_ _01219_ _01438_ _01842_ VGND VGND VPWR VPWR _01853_ sky130_fd_sc_hd__or4_4
XFILLER_0_116_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07809__D _06637_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_711 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07158_ _01065_ _01087_ VGND VGND VPWR VPWR _01098_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_89_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07089_ _00333_ VGND VGND VPWR VPWR _00344_ sky130_fd_sc_hd__buf_6
XANTENNA__07394__A net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10251__C _02482_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09106__A1 _00530_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12810_ _05108_ _05114_ _05099_ VGND VGND VPWR VPWR _05296_ sky130_fd_sc_hd__o21a_1
XANTENNA__07841__B _06967_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13790_ _06331_ _06355_ VGND VGND VPWR VPWR _06356_ sky130_fd_sc_hd__and2_1
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12741_ _00783_ _00779_ _02133_ VGND VGND VPWR VPWR _05220_ sky130_fd_sc_hd__and3_1
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12672_ _05119_ _05143_ VGND VGND VPWR VPWR _05144_ sky130_fd_sc_hd__xnor2_1
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08953__A _01061_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11623_ _03987_ _03989_ VGND VGND VPWR VPWR _03990_ sky130_fd_sc_hd__nand2_1
XTAP_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07569__A _01361_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11554_ _03510_ _06874_ _01177_ VGND VGND VPWR VPWR _03914_ sky130_fd_sc_hd__and3_1
XFILLER_0_108_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10505_ _02760_ VGND VGND VPWR VPWR _02761_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11485_ _03811_ _03836_ _03837_ VGND VGND VPWR VPWR _03838_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_123_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_711 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13224_ _05648_ _05747_ _05750_ VGND VGND VPWR VPWR _05751_ sky130_fd_sc_hd__a21o_1
XFILLER_0_122_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10436_ _02684_ _02685_ VGND VGND VPWR VPWR _02687_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11819__A _00157_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09593__A1 _03685_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13155_ _05668_ _05671_ _05674_ VGND VGND VPWR VPWR _05675_ sky130_fd_sc_hd__a21o_1
X_10367_ _02608_ _02610_ VGND VGND VPWR VPWR _02611_ sky130_fd_sc_hd__nand2_1
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12106_ _03997_ _04520_ VGND VGND VPWR VPWR _04522_ sky130_fd_sc_hd__nor2_2
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10298_ _02329_ _02533_ VGND VGND VPWR VPWR _02535_ sky130_fd_sc_hd__or2_1
X_13086_ _05474_ _05490_ VGND VGND VPWR VPWR _05600_ sky130_fd_sc_hd__or2_1
X_12037_ _04382_ _04383_ _04384_ _04380_ VGND VGND VPWR VPWR _04446_ sky130_fd_sc_hd__a31o_1
XANTENNA__07454__D _02982_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11554__A _03510_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13988_ _06565_ _06569_ VGND VGND VPWR VPWR _06574_ sky130_fd_sc_hd__nor2_1
XFILLER_0_125_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09024__A _03543_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12939_ _04566_ _04583_ _04574_ VGND VGND VPWR VPWR _05438_ sky130_fd_sc_hd__or3_1
XFILLER_0_48_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08130_ _07039_ _07075_ _00077_ _00173_ VGND VGND VPWR VPWR _00174_ sky130_fd_sc_hd__a31o_2
XFILLER_0_44_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08061_ _05588_ _06744_ _00103_ _00104_ VGND VGND VPWR VPWR _00105_ sky130_fd_sc_hd__and4_1
XFILLER_0_113_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08387__A2 _00373_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08963_ _04169_ _01076_ net47 net48 VGND VGND VPWR VPWR _01073_ sky130_fd_sc_hd__and4_1
XANTENNA__11448__B _03683_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07914_ _00901_ _04455_ _06917_ VGND VGND VPWR VPWR _07043_ sky130_fd_sc_hd__and3_1
X_08894_ _00807_ _00809_ _00508_ _00298_ VGND VGND VPWR VPWR _00998_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_75_61 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12340__B1 _00959_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07845_ _06872_ _06880_ _06864_ VGND VGND VPWR VPWR _06974_ sky130_fd_sc_hd__a21o_1
XFILLER_0_75_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11464__A _00497_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07776_ net33 net6 _05005_ _04994_ VGND VGND VPWR VPWR _06905_ sky130_fd_sc_hd__a31o_1
XFILLER_0_78_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09639__A2 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09515_ _01535_ _01676_ VGND VGND VPWR VPWR _01677_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11446__A2 _03682_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_736 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09869__A _06964_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09446_ _02335_ _01601_ VGND VGND VPWR VPWR _01603_ sky130_fd_sc_hd__nand2_1
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11911__B _06450_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09377_ _01501_ _01526_ VGND VGND VPWR VPWR _01527_ sky130_fd_sc_hd__nor2_1
XANTENNA__12295__A _02188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08328_ _00379_ VGND VGND VPWR VPWR _00380_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_117_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10957__A1 _00145_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08259_ _06417_ _00138_ _04906_ _04928_ VGND VGND VPWR VPWR _00304_ sky130_fd_sc_hd__and4_1
XFILLER_0_104_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11270_ _03591_ _03592_ VGND VGND VPWR VPWR _03603_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_120_705 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10221_ _02029_ _01564_ _02449_ _02450_ VGND VGND VPWR VPWR _02451_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_30_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10543__A _00388_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_574 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10185__A2 net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10152_ _02364_ _02374_ VGND VGND VPWR VPWR _02375_ sky130_fd_sc_hd__xnor2_4
X_10083_ _02236_ _02239_ VGND VGND VPWR VPWR _02299_ sky130_fd_sc_hd__or2b_1
XANTENNA__08948__A _00410_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13911_ _06234_ _06201_ _06231_ VGND VGND VPWR VPWR _06489_ sky130_fd_sc_hd__or3_1
XANTENNA__11374__A _01312_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13842_ _06376_ _06412_ VGND VGND VPWR VPWR _06413_ sky130_fd_sc_hd__nor2_1
XFILLER_0_69_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12634__A1 _02168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13773_ _06268_ _06336_ VGND VGND VPWR VPWR _06337_ sky130_fd_sc_hd__or2_1
X_10985_ _03278_ _03288_ VGND VGND VPWR VPWR _03289_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_427 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12724_ _05199_ _05200_ VGND VGND VPWR VPWR _05201_ sky130_fd_sc_hd__or2b_1
XANTENNA__09779__A _01197_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08683__A _00563_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12655_ _05119_ _05123_ _05124_ VGND VGND VPWR VPWR _05125_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_127_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11606_ _03970_ _03964_ VGND VGND VPWR VPWR _03972_ sky130_fd_sc_hd__nor2_1
X_12586_ _03707_ _03740_ _02158_ _02304_ VGND VGND VPWR VPWR _05050_ sky130_fd_sc_hd__and4_1
XFILLER_0_37_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11537_ _06873_ _01178_ _01247_ _06874_ VGND VGND VPWR VPWR _03896_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_41_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_output97_A net97 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11468_ _00497_ _02673_ VGND VGND VPWR VPWR _03820_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap139 net180 VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__buf_1
XANTENNA__12652__B _02759_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08369__A2 _00423_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13207_ _05725_ _05732_ VGND VGND VPWR VPWR _05733_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10419_ _01295_ net21 _02133_ _01306_ VGND VGND VPWR VPWR _02668_ sky130_fd_sc_hd__a22o_1
X_14187_ _06627_ _06786_ VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__xnor2_4
XFILLER_0_21_574 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11399_ _02120_ VGND VGND VPWR VPWR _03744_ sky130_fd_sc_hd__clkbuf_4
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09019__A _06965_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13138_ _05209_ _05210_ _05656_ VGND VGND VPWR VPWR _05657_ sky130_fd_sc_hd__a21oi_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13069_ _05563_ _05580_ VGND VGND VPWR VPWR _05581_ sky130_fd_sc_hd__nand2_1
XANTENNA__08858__A net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07630_ _06186_ _06252_ VGND VGND VPWR VPWR _06263_ sky130_fd_sc_hd__and2_1
XFILLER_0_45_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07481__B _04598_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07561_ _05511_ _05423_ VGND VGND VPWR VPWR _05522_ sky130_fd_sc_hd__and2b_1
XANTENNA__12625__A1 _00572_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12625__B2 _00414_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09300_ _01170_ _01171_ _01440_ VGND VGND VPWR VPWR _01442_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_75_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07492_ _04741_ _04752_ VGND VGND VPWR VPWR _04763_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_146_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09231_ _01339_ _00604_ _01074_ _01073_ VGND VGND VPWR VPWR _01367_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_118_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09460__A1_N _00475_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12389__B1 _01584_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09201__B _06966_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09162_ _03070_ _02280_ _00416_ _01288_ VGND VGND VPWR VPWR _01291_ sky130_fd_sc_hd__and4_1
XFILLER_0_71_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08113_ _01361_ VGND VGND VPWR VPWR _00157_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_44_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09093_ _01206_ _01215_ VGND VGND VPWR VPWR _01216_ sky130_fd_sc_hd__xor2_1
XFILLER_0_31_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07359__D _02719_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08044_ _07079_ _07080_ _07001_ VGND VGND VPWR VPWR _00088_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_31_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10363__A _06744_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09995_ _01904_ _02202_ VGND VGND VPWR VPWR _02203_ sky130_fd_sc_hd__or2_1
X_08946_ _00898_ _01054_ VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__xor2_2
X_08877_ _00775_ _00977_ _00979_ VGND VGND VPWR VPWR _00980_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_99_828 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07828_ _00880_ net36 _06866_ _06865_ VGND VGND VPWR VPWR _06957_ sky130_fd_sc_hd__a31o_1
X_07759_ _00453_ _06885_ _06887_ VGND VGND VPWR VPWR _06888_ sky130_fd_sc_hd__nand3_1
XFILLER_0_39_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10770_ _02933_ _03052_ VGND VGND VPWR VPWR _03053_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_137_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09429_ _01211_ VGND VGND VPWR VPWR _01584_ sky130_fd_sc_hd__buf_4
XFILLER_0_94_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08048__A1 _03521_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12440_ _04769_ _04888_ VGND VGND VPWR VPWR _04889_ sky130_fd_sc_hd__nand2_1
XANTENNA__08048__B2 _00377_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_817 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12371_ _04803_ _04802_ VGND VGND VPWR VPWR _04813_ sky130_fd_sc_hd__and2b_1
XFILLER_0_133_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12753__A _01507_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14110_ _06077_ _04013_ VGND VGND VPWR VPWR _06706_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11322_ _02933_ _03052_ _03659_ VGND VGND VPWR VPWR _03660_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_120_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14041_ _06630_ _06631_ VGND VGND VPWR VPWR _06632_ sky130_fd_sc_hd__nand2_4
XFILLER_0_31_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11253_ _03578_ _03582_ _03583_ VGND VGND VPWR VPWR _03584_ sky130_fd_sc_hd__or3_1
XANTENNA__10273__A _03576_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10204_ _02425_ _02101_ _02430_ VGND VGND VPWR VPWR _02432_ sky130_fd_sc_hd__o21a_1
X_11184_ _03041_ _03507_ VGND VGND VPWR VPWR _03508_ sky130_fd_sc_hd__nor2_1
X_10135_ _02971_ net46 _01368_ _00366_ VGND VGND VPWR VPWR _02356_ sky130_fd_sc_hd__a22o_1
XANTENNA__09781__B net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07582__A _05731_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10066_ _01752_ _01867_ VGND VGND VPWR VPWR _02281_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10330__A2 net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13825_ _06379_ _06393_ VGND VGND VPWR VPWR _06394_ sky130_fd_sc_hd__or2_1
XANTENNA__13804__B1 _03680_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13756_ _06305_ _06317_ VGND VGND VPWR VPWR _06319_ sky130_fd_sc_hd__nor2_1
X_10968_ _04862_ net4 net46 _01368_ VGND VGND VPWR VPWR _03271_ sky130_fd_sc_hd__and4_1
XFILLER_0_73_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12707_ _05077_ VGND VGND VPWR VPWR _05183_ sky130_fd_sc_hd__inv_2
X_13687_ _01288_ _02090_ _02725_ _02728_ VGND VGND VPWR VPWR _06243_ sky130_fd_sc_hd__and4_1
XFILLER_0_128_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10899_ _03163_ _03159_ _03161_ VGND VGND VPWR VPWR _03195_ sky130_fd_sc_hd__nor3_1
XFILLER_0_5_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09021__B _06966_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12638_ _05105_ _05040_ VGND VGND VPWR VPWR _05107_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13583__A2 _02858_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12569_ _05003_ _05029_ _05030_ VGND VGND VPWR VPWR _05031_ sky130_fd_sc_hd__a21o_1
XFILLER_0_13_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13335__A2 _02724_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08800_ _00895_ _00569_ _00720_ _00566_ VGND VGND VPWR VPWR _00896_ sky130_fd_sc_hd__a211o_2
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09691__B _04059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09780_ _01965_ _01966_ _01967_ VGND VGND VPWR VPWR _01968_ sky130_fd_sc_hd__a21oi_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08731_ _00263_ _00819_ VGND VGND VPWR VPWR _00820_ sky130_fd_sc_hd__nand2_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10630__B _02731_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09711__A1 _06461_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08662_ _00157_ _00741_ _00743_ _00583_ VGND VGND VPWR VPWR _00744_ sky130_fd_sc_hd__and4_1
XANTENNA__11445__C _03682_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07613_ net187 _05988_ _06054_ VGND VGND VPWR VPWR _06076_ sky130_fd_sc_hd__nand3_4
X_08593_ _06494_ _00004_ _00471_ _00472_ VGND VGND VPWR VPWR _00669_ sky130_fd_sc_hd__a31o_1
XFILLER_0_49_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07544_ _05324_ _04796_ VGND VGND VPWR VPWR _05335_ sky130_fd_sc_hd__xnor2_2
XANTENNA__13271__A1 _05773_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_717 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11461__B _00121_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07475_ _04411_ _04477_ _04554_ VGND VGND VPWR VPWR _04576_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_119_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09214_ _01316_ _01347_ VGND VGND VPWR VPWR _01348_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_91_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09145_ net15 VGND VGND VPWR VPWR _01272_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_16_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09076_ _01996_ net11 _01194_ _01195_ VGND VGND VPWR VPWR _01198_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_130_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08027_ _00069_ _00070_ VGND VGND VPWR VPWR _00071_ sky130_fd_sc_hd__and2_1
XFILLER_0_141_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07386__B _03587_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09978_ _01891_ _01898_ VGND VGND VPWR VPWR _02185_ sky130_fd_sc_hd__or2b_1
XANTENNA__07961__B1 _07004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08929_ _00866_ VGND VGND VPWR VPWR _01037_ sky130_fd_sc_hd__inv_2
XANTENNA__10540__B _02169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10848__B1 net52 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11940_ _04337_ _04338_ VGND VGND VPWR VPWR _04339_ sky130_fd_sc_hd__nor2_1
XANTENNA__11355__C _01312_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11871_ _00004_ _01601_ _04258_ _04259_ VGND VGND VPWR VPWR _04263_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_95_820 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13610_ _06138_ _06148_ _06149_ _06147_ VGND VGND VPWR VPWR _06158_ sky130_fd_sc_hd__o22a_1
X_10822_ _03587_ _00891_ net56 net57 VGND VGND VPWR VPWR _03110_ sky130_fd_sc_hd__and4_1
XFILLER_0_79_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13541_ _06048_ _06073_ _06081_ VGND VGND VPWR VPWR _06082_ sky130_fd_sc_hd__a21oi_1
X_10753_ _00399_ _02765_ _03033_ VGND VGND VPWR VPWR _03034_ sky130_fd_sc_hd__a21o_1
XFILLER_0_137_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13472_ _05993_ _05989_ _06004_ VGND VGND VPWR VPWR _06006_ sky130_fd_sc_hd__and3_1
XFILLER_0_54_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10684_ _02945_ _02957_ VGND VGND VPWR VPWR _02958_ sky130_fd_sc_hd__nor2_1
XFILLER_0_109_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12423_ _04858_ _04859_ _04869_ VGND VGND VPWR VPWR _04870_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_35_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12483__A _00612_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10379__A2 _00734_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08441__A1 _03059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12354_ _04790_ _04793_ VGND VGND VPWR VPWR _04794_ sky130_fd_sc_hd__and2b_1
XANTENNA__09495__C net50 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11305_ _03634_ _03636_ VGND VGND VPWR VPWR _03641_ sky130_fd_sc_hd__nor2_1
X_12285_ _04714_ _01181_ _04716_ VGND VGND VPWR VPWR _04718_ sky130_fd_sc_hd__and3_1
X_14024_ _05750_ _06611_ _06612_ VGND VGND VPWR VPWR _06613_ sky130_fd_sc_hd__a21o_1
X_11236_ _02979_ _03564_ VGND VGND VPWR VPWR _03566_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11167_ _03468_ _03487_ _03489_ VGND VGND VPWR VPWR _03490_ sky130_fd_sc_hd__o21a_1
X_10118_ _06637_ _02190_ _02337_ VGND VGND VPWR VPWR _02338_ sky130_fd_sc_hd__and3_1
XFILLER_0_93_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11098_ _01400_ VGND VGND VPWR VPWR _03414_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__13464__D _02731_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10049_ _01855_ _02262_ VGND VGND VPWR VPWR _02263_ sky130_fd_sc_hd__nand2_1
XFILLER_0_117_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13808_ _06374_ _06375_ VGND VGND VPWR VPWR _06376_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09457__B1 net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13739_ _05858_ _06297_ _06299_ VGND VGND VPWR VPWR _06300_ sky130_fd_sc_hd__and3_1
XFILLER_0_46_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09967__A _01934_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07260_ _02094_ _02193_ _02204_ VGND VGND VPWR VPWR _02215_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_73_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07191_ _01251_ _01241_ VGND VGND VPWR VPWR _01459_ sky130_fd_sc_hd__or2b_4
XFILLER_0_143_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09901_ _02098_ _02099_ VGND VGND VPWR VPWR _02100_ sky130_fd_sc_hd__nor2_1
XFILLER_0_111_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09832_ _07004_ _00390_ _02024_ VGND VGND VPWR VPWR _02025_ sky130_fd_sc_hd__and3_1
XANTENNA__11417__A1_N _00003_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10542__A2 _02724_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09763_ _01716_ _01717_ _01945_ VGND VGND VPWR VPWR _01949_ sky130_fd_sc_hd__and3_2
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10360__B _03773_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08714_ _00775_ _00800_ VGND VGND VPWR VPWR _00801_ sky130_fd_sc_hd__xnor2_1
X_09694_ _04378_ _04103_ _00777_ _02971_ VGND VGND VPWR VPWR _01873_ sky130_fd_sc_hd__a22oi_1
Xrebuffer10 _01799_ VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrebuffer21 net183 VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer32 _06065_ VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_96_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08645_ _00725_ VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07171__A1 _00978_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07171__B2 _00869_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08576_ _00648_ _00649_ VGND VGND VPWR VPWR _00651_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07527_ _04345_ _05115_ _05137_ VGND VGND VPWR VPWR _05148_ sky130_fd_sc_hd__or3_4
XFILLER_0_76_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10088__A _02304_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_763 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07458_ net58 net31 net32 net175 VGND VGND VPWR VPWR _04389_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_344 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_638 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07389_ _03048_ _03620_ VGND VGND VPWR VPWR _03631_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_17_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10816__A _06637_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__07397__A net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09128_ _01247_ VGND VGND VPWR VPWR _01254_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_32_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09059_ _01178_ VGND VGND VPWR VPWR _01179_ sky130_fd_sc_hd__buf_4
XFILLER_0_60_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12070_ _04465_ _04474_ _04478_ VGND VGND VPWR VPWR _04482_ sky130_fd_sc_hd__and3_1
XANTENNA__11647__A _02246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11021_ _03316_ _03319_ _03320_ VGND VGND VPWR VPWR _03329_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11191__C1 _01108_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12972_ _05451_ _05473_ VGND VGND VPWR VPWR _05474_ sky130_fd_sc_hd__xnor2_4
XANTENNA__08956__A _00460_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12286__A2 _01956_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11923_ _04318_ _04319_ VGND VGND VPWR VPWR _04320_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11382__A _02246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11854_ _04234_ _04243_ VGND VGND VPWR VPWR _04244_ sky130_fd_sc_hd__xor2_1
XFILLER_0_68_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10805_ _03089_ _03090_ VGND VGND VPWR VPWR _03091_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11785_ _04165_ _02657_ _04166_ VGND VGND VPWR VPWR _04168_ sky130_fd_sc_hd__a21o_1
XFILLER_0_55_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13524_ _06060_ _06061_ _06036_ _06037_ VGND VGND VPWR VPWR _06063_ sky130_fd_sc_hd__a211oi_1
XANTENNA__12994__B1 _00381_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10736_ _03006_ _03011_ _03014_ VGND VGND VPWR VPWR _03016_ sky130_fd_sc_hd__and3_1
XFILLER_0_94_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13455_ _05984_ _05986_ VGND VGND VPWR VPWR _05987_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_82_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10667_ _05192_ _01546_ _02156_ _02982_ VGND VGND VPWR VPWR _02940_ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_479 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12406_ _00782_ _00413_ _00571_ _00373_ VGND VGND VPWR VPWR _04852_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13386_ _05910_ _05911_ VGND VGND VPWR VPWR _05913_ sky130_fd_sc_hd__nor2_1
X_10598_ _02862_ _02863_ VGND VGND VPWR VPWR _02864_ sky130_fd_sc_hd__nor2_1
XFILLER_0_112_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07100__A _00453_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput108 net108 VGND VGND VPWR VPWR prod[49] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12337_ _04771_ _04770_ VGND VGND VPWR VPWR _04776_ sky130_fd_sc_hd__and2b_1
XFILLER_0_23_488 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput119 net119 VGND VGND VPWR VPWR prod[59] sky130_fd_sc_hd__buf_6
XANTENNA__10772__A2 _02724_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12268_ _04649_ _04699_ VGND VGND VPWR VPWR _04700_ sky130_fd_sc_hd__xor2_1
XFILLER_0_120_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14007_ _06594_ VGND VGND VPWR VPWR _06595_ sky130_fd_sc_hd__inv_2
X_11219_ _00410_ _01108_ VGND VGND VPWR VPWR _03547_ sky130_fd_sc_hd__nand2_2
X_12199_ _04610_ _04613_ _04618_ _04623_ VGND VGND VPWR VPWR _04624_ sky130_fd_sc_hd__o211ai_4
Xoutput90 net90 VGND VGND VPWR VPWR prod[32] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_78_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12388__A _00784_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08430_ _00487_ _00489_ VGND VGND VPWR VPWR _00491_ sky130_fd_sc_hd__and2_1
XFILLER_0_53_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08361_ _00414_ VGND VGND VPWR VPWR _00415_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_18_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__11788__A1 _02127_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07312_ _02762_ _02773_ VGND VGND VPWR VPWR _02784_ sky130_fd_sc_hd__and2b_1
XANTENNA__11788__B2 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09697__A _04598_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08292_ _00098_ _00339_ VGND VGND VPWR VPWR _00340_ sky130_fd_sc_hd__nand2_2
XFILLER_0_74_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12835__B _01933_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07243_ _00901_ VGND VGND VPWR VPWR _02029_ sky130_fd_sc_hd__buf_4
XFILLER_0_144_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_254 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07174_ _01219_ VGND VGND VPWR VPWR _01273_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09090__A2_N _01211_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_140 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13701__A2 _02721_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09815_ _02003_ _02005_ VGND VGND VPWR VPWR _02006_ sky130_fd_sc_hd__xor2_2
XANTENNA__10090__B _02306_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09746_ _01928_ _01929_ VGND VGND VPWR VPWR _01931_ sky130_fd_sc_hd__or2b_1
XANTENNA__09133__A2 _03773_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09677_ _01838_ _01854_ VGND VGND VPWR VPWR _01855_ sky130_fd_sc_hd__and2_1
XTAP_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07144__A1 _00420_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08341__B1 _00393_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08628_ _00466_ _00524_ _00547_ VGND VGND VPWR VPWR _00708_ sky130_fd_sc_hd__a21o_1
XFILLER_0_96_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08559_ _00410_ _00544_ _00542_ VGND VGND VPWR VPWR _00632_ sky130_fd_sc_hd__nand3_1
XTAP_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11570_ _03930_ _03931_ VGND VGND VPWR VPWR _03932_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10521_ _02777_ _02778_ VGND VGND VPWR VPWR _02779_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13240_ _05762_ _05764_ _05765_ VGND VGND VPWR VPWR _05766_ sky130_fd_sc_hd__and3_1
XFILLER_0_107_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10452_ _02592_ _02593_ _02703_ VGND VGND VPWR VPWR _02704_ sky130_fd_sc_hd__nand3_1
XANTENNA__08016__A _01197_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13171_ _05690_ _05691_ _05692_ VGND VGND VPWR VPWR _05693_ sky130_fd_sc_hd__a21o_2
XFILLER_0_103_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10383_ _02623_ _02626_ VGND VGND VPWR VPWR _02628_ sky130_fd_sc_hd__or2_1
XFILLER_0_103_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12122_ _04002_ _04538_ VGND VGND VPWR VPWR _04539_ sky130_fd_sc_hd__nor2_1
XFILLER_0_102_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13576__B _03785_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12053_ _04247_ _04249_ _04244_ VGND VGND VPWR VPWR _04463_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10506__A2 _02721_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11004_ _04598_ _01506_ _01369_ _05203_ VGND VGND VPWR VPWR _03310_ sky130_fd_sc_hd__a22oi_1
XANTENNA__07383__A1 _00453_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07383__B2 _02051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08580__B1 _00543_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08686__A _05577_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12955_ _05454_ _05029_ VGND VGND VPWR VPWR _05455_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_99_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11906_ _04299_ _04300_ VGND VGND VPWR VPWR _04302_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12886_ _05377_ _05378_ VGND VGND VPWR VPWR _05380_ sky130_fd_sc_hd__and2_1
XTAP_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11837_ _04193_ _04225_ VGND VGND VPWR VPWR _04226_ sky130_fd_sc_hd__and2_1
XTAP_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11768_ _04148_ _04149_ VGND VGND VPWR VPWR _04150_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_56_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13507_ _06025_ _06028_ _06042_ VGND VGND VPWR VPWR _06045_ sky130_fd_sc_hd__and3_1
X_10719_ _02924_ _02996_ VGND VGND VPWR VPWR _02997_ sky130_fd_sc_hd__and2_1
XFILLER_0_130_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11699_ _04072_ _04073_ VGND VGND VPWR VPWR _04074_ sky130_fd_sc_hd__nor2_1
XANTENNA__12374__C _00457_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13438_ _03785_ VGND VGND VPWR VPWR _05969_ sky130_fd_sc_hd__buf_2
XANTENNA__08571__D _00151_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xrebuffer1 _03235_ VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_113_416 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07468__C _04378_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_252 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13369_ _05892_ _05893_ VGND VGND VPWR VPWR _05894_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_279 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07930_ net163 net6 net5 _00705_ VGND VGND VPWR VPWR _07059_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_48_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09980__A _01664_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07861_ _06142_ _06175_ _06406_ VGND VGND VPWR VPWR _06990_ sky130_fd_sc_hd__a21oi_1
X_09600_ _01302_ _01620_ _01770_ VGND VGND VPWR VPWR _01771_ sky130_fd_sc_hd__nor3_1
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07792_ _05148_ _06920_ VGND VGND VPWR VPWR _06921_ sky130_fd_sc_hd__nor2_2
XANTENNA__08596__A _06472_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09531_ _01541_ _01543_ _01694_ VGND VGND VPWR VPWR _01695_ sky130_fd_sc_hd__a21o_1
XANTENNA__07931__C net6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09462_ _01618_ _01619_ VGND VGND VPWR VPWR _01620_ sky130_fd_sc_hd__or2_2
XANTENNA__11453__C _03532_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08413_ _02149_ _05577_ _07010_ _00101_ VGND VGND VPWR VPWR _00472_ sky130_fd_sc_hd__and4_1
XFILLER_0_19_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10681__A1 _00094_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09393_ _01541_ _01543_ VGND VGND VPWR VPWR _01544_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_46_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08344_ _00354_ _00368_ VGND VGND VPWR VPWR _00397_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_74_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11630__B1 _01155_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08275_ _00319_ _00320_ VGND VGND VPWR VPWR _00321_ sky130_fd_sc_hd__and2_1
XFILLER_0_73_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07226_ _01448_ _01832_ VGND VGND VPWR VPWR _01842_ sky130_fd_sc_hd__and2_4
XFILLER_0_116_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_736 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07157_ _01076_ net60 VGND VGND VPWR VPWR _01087_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11933__A1 _00113_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07675__A _00442_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07088_ _00322_ VGND VGND VPWR VPWR _00333_ sky130_fd_sc_hd__buf_4
XANTENNA__09890__A _01780_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09106__A2 _00391_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09729_ _01910_ _01911_ VGND VGND VPWR VPWR _01912_ sky130_fd_sc_hd__nor2_2
XANTENNA__13562__D _02736_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12740_ _04633_ _04635_ _04637_ VGND VGND VPWR VPWR _05219_ sky130_fd_sc_hd__or3b_1
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12671_ _05124_ _05123_ VGND VGND VPWR VPWR _05143_ sky130_fd_sc_hd__nand2_1
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12756__A _00607_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11622_ _00519_ _01957_ _03988_ VGND VGND VPWR VPWR _03989_ sky130_fd_sc_hd__a21o_1
XTAP_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11553_ _06874_ _01177_ _01247_ _03510_ VGND VGND VPWR VPWR _03913_ sky130_fd_sc_hd__a22o_1
XANTENNA__10276__A _04081_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07569__B _05566_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10504_ _00635_ _07040_ _02720_ _02726_ VGND VGND VPWR VPWR _02760_ sky130_fd_sc_hd__and4_1
X_11484_ _03797_ _03799_ VGND VGND VPWR VPWR _03837_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13223_ _05628_ _05630_ _05749_ VGND VGND VPWR VPWR _05750_ sky130_fd_sc_hd__o21a_1
X_10435_ _02447_ _02457_ _02469_ VGND VGND VPWR VPWR _02685_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_21_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13154_ _05208_ _05673_ VGND VGND VPWR VPWR _05674_ sky130_fd_sc_hd__xnor2_4
XANTENNA__11819__B _03678_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10366_ _02604_ _02607_ VGND VGND VPWR VPWR _02610_ sky130_fd_sc_hd__or2_1
X_12105_ _03996_ _03983_ _03994_ VGND VGND VPWR VPWR _04520_ sky130_fd_sc_hd__and3_1
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13085_ _05453_ _05471_ VGND VGND VPWR VPWR _05598_ sky130_fd_sc_hd__nand2_1
X_10297_ _02329_ _02533_ VGND VGND VPWR VPWR _02534_ sky130_fd_sc_hd__nand2_1
XANTENNA__11538__C _03510_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12036_ _04442_ _04443_ VGND VGND VPWR VPWR _04445_ sky130_fd_sc_hd__nand2_1
XANTENNA__14211__A _06800_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11554__B _06874_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13987_ _05946_ _06563_ _06572_ VGND VGND VPWR VPWR _06573_ sky130_fd_sc_hd__o21a_1
XANTENNA__09024__B _00298_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12938_ _04570_ _04571_ _02473_ _02475_ _02699_ VGND VGND VPWR VPWR _05437_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_125_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12869_ _05320_ _05321_ _05359_ VGND VGND VPWR VPWR _05361_ sky130_fd_sc_hd__nand3_1
XFILLER_0_145_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_344 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11612__B1 _03687_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07479__B net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08060_ _02105_ _00101_ _06733_ _00650_ VGND VGND VPWR VPWR _00104_ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_780 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07595__A1 _02029_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08962_ _04081_ _00604_ _00960_ _00958_ VGND VGND VPWR VPWR _01072_ sky130_fd_sc_hd__a31o_1
X_07913_ _06911_ _06927_ VGND VGND VPWR VPWR _07042_ sky130_fd_sc_hd__nand2_1
X_08893_ _00995_ _00996_ VGND VGND VPWR VPWR _00997_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12340__A1 _03762_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07844_ _06951_ _06972_ VGND VGND VPWR VPWR _06973_ sky130_fd_sc_hd__xor2_1
XFILLER_0_75_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11464__B _03681_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07775_ _06902_ _06903_ VGND VGND VPWR VPWR _06904_ sky130_fd_sc_hd__xnor2_1
X_09514_ _01674_ _01675_ VGND VGND VPWR VPWR _01676_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09445_ _01600_ VGND VGND VPWR VPWR _01601_ sky130_fd_sc_hd__clkbuf_4
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09869__B _00121_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09376_ _01515_ _01524_ VGND VGND VPWR VPWR _01526_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11911__C _03750_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12295__B _02427_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10406__A1 _02029_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08327_ _00378_ VGND VGND VPWR VPWR _00379_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_117_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10957__A2 _00608_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08258_ _00291_ _00302_ VGND VGND VPWR VPWR _00303_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07209_ _01635_ _01645_ VGND VGND VPWR VPWR _01656_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10824__A _01372_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08189_ _00224_ _00231_ _00232_ VGND VGND VPWR VPWR _00233_ sky130_fd_sc_hd__a21o_2
XFILLER_0_104_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10220_ _05467_ _01000_ _01177_ _01246_ VGND VGND VPWR VPWR _02450_ sky130_fd_sc_hd__and4_1
XFILLER_0_120_739 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10543__B _03004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10151_ _02372_ _02373_ VGND VGND VPWR VPWR _02374_ sky130_fd_sc_hd__nor2_2
XANTENNA__09109__B _01233_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10082_ _00991_ _01356_ _01756_ _01757_ _02297_ VGND VGND VPWR VPWR _02298_ sky130_fd_sc_hd__a311o_1
XANTENNA__08948__B _00380_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13910_ net137 net136 VGND VGND VPWR VPWR _06488_ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11374__B _00544_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09125__A _01249_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13841_ _06374_ _06375_ VGND VGND VPWR VPWR _06412_ sky130_fd_sc_hd__nor2_1
XFILLER_0_69_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13772_ _02765_ _05887_ _06267_ VGND VGND VPWR VPWR _06336_ sky130_fd_sc_hd__a21oi_1
X_10984_ _03286_ _03287_ VGND VGND VPWR VPWR _03288_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12723_ _00391_ _01062_ _05197_ VGND VGND VPWR VPWR _05200_ sky130_fd_sc_hd__a21o_1
XANTENNA__09779__B _04510_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08683__B _00639_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_316 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12654_ _00390_ _02759_ _05121_ VGND VGND VPWR VPWR _05124_ sky130_fd_sc_hd__a21o_1
XFILLER_0_38_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11605_ _03967_ VGND VGND VPWR VPWR _03970_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09263__A1 _01066_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12585_ _03740_ _02158_ _02304_ _03707_ VGND VGND VPWR VPWR _05048_ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11540__D net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09795__A _05456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11536_ _06819_ _06874_ _01177_ _01247_ VGND VGND VPWR VPWR _03895_ sky130_fd_sc_hd__and4_1
XFILLER_0_135_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11467_ _03803_ _03818_ VGND VGND VPWR VPWR _03819_ sky130_fd_sc_hd__or2_1
X_13206_ _05728_ _05730_ VGND VGND VPWR VPWR _05732_ sky130_fd_sc_hd__xor2_2
XFILLER_0_110_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10418_ _01295_ _01306_ net22 VGND VGND VPWR VPWR _02667_ sky130_fd_sc_hd__and3_1
X_14186_ _06623_ _06643_ _06757_ _06784_ _05968_ VGND VGND VPWR VPWR _06786_ sky130_fd_sc_hd__o32a_2
X_11398_ _03741_ _03742_ VGND VGND VPWR VPWR _03743_ sky130_fd_sc_hd__and2b_1
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_586 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13137_ _05182_ _05208_ _05211_ VGND VGND VPWR VPWR _05656_ sky130_fd_sc_hd__o21a_1
X_10349_ _02589_ _02590_ VGND VGND VPWR VPWR _02591_ sky130_fd_sc_hd__nand2_1
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09019__B _04906_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13068_ _05575_ _05579_ VGND VGND VPWR VPWR _05580_ sky130_fd_sc_hd__and2_1
X_12019_ _04353_ _04354_ _04355_ _04351_ VGND VGND VPWR VPWR _04426_ sky130_fd_sc_hd__a31o_1
XANTENNA__11565__A _00486_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07560_ _05434_ _05500_ VGND VGND VPWR VPWR _05511_ sky130_fd_sc_hd__xor2_2
XANTENNA__12625__A2 _01411_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09689__B _01867_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07491_ _04620_ _04609_ VGND VGND VPWR VPWR _04752_ sky130_fd_sc_hd__and2b_1
XFILLER_0_88_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09230_ _01071_ _01079_ VGND VGND VPWR VPWR _01366_ sky130_fd_sc_hd__and2b_1
XFILLER_0_146_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12389__A1 _00779_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09161_ _03070_ _01188_ _01289_ _02456_ VGND VGND VPWR VPWR _01290_ sky130_fd_sc_hd__a22o_1
XANTENNA__12389__B2 _00784_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09201__C _00143_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08112_ _00154_ _00155_ VGND VGND VPWR VPWR _00156_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_126_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09092_ _01207_ _01214_ VGND VGND VPWR VPWR _01215_ sky130_fd_sc_hd__xor2_1
XFILLER_0_114_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08043_ _07079_ _07080_ VGND VGND VPWR VPWR _00087_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08114__A net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10363__B _03938_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09994_ _02200_ _02201_ VGND VGND VPWR VPWR _02202_ sky130_fd_sc_hd__nor2_1
XFILLER_0_110_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08945_ _00899_ _01053_ VGND VGND VPWR VPWR _01054_ sky130_fd_sc_hd__xnor2_4
XANTENNA__12313__A1 _00459_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12313__B2 _01288_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08876_ _00789_ _00799_ VGND VGND VPWR VPWR _00979_ sky130_fd_sc_hd__nand2_1
X_07827_ _06954_ _06955_ VGND VGND VPWR VPWR _06956_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07758_ _06886_ _06847_ VGND VGND VPWR VPWR _06887_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13813__A1 _03414_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07689_ net35 VGND VGND VPWR VPWR _06818_ sky130_fd_sc_hd__clkbuf_4
X_09428_ _01207_ _01214_ _01278_ VGND VGND VPWR VPWR _01583_ sky130_fd_sc_hd__and3_1
XFILLER_0_94_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09359_ _01506_ VGND VGND VPWR VPWR _01507_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_34_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09245__A1 _05566_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08048__A2 _02993_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12370_ _04809_ _04810_ VGND VGND VPWR VPWR _04812_ sky130_fd_sc_hd__xor2_1
XFILLER_0_105_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12753__B _01504_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11321_ _02920_ _02932_ VGND VGND VPWR VPWR _03659_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14040_ net135 _06578_ _06629_ VGND VGND VPWR VPWR _06631_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_132_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11252_ _03545_ _03581_ _03580_ VGND VGND VPWR VPWR _03583_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10273__B _00989_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10203_ _02425_ _02101_ _02430_ VGND VGND VPWR VPWR _02431_ sky130_fd_sc_hd__nor3_1
X_11183_ _03038_ _03040_ VGND VGND VPWR VPWR _03507_ sky130_fd_sc_hd__and2_1
X_10134_ _02353_ _02354_ VGND VGND VPWR VPWR _02355_ sky130_fd_sc_hd__xnor2_2
XANTENNA__08508__B1 _00575_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07582__B _01000_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10065_ _02055_ _02272_ VGND VGND VPWR VPWR _02279_ sky130_fd_sc_hd__nor2_2
XFILLER_0_106_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13824_ _03414_ _03683_ _06377_ _06378_ VGND VGND VPWR VPWR _06393_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__12068__B1 _01252_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13804__A1 _02190_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08694__A _00778_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13804__B2 _02188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10967_ _03260_ _03267_ VGND VGND VPWR VPWR _03270_ sky130_fd_sc_hd__xor2_1
X_13755_ _05875_ _05881_ _06304_ VGND VGND VPWR VPWR _06317_ sky130_fd_sc_hd__nor3_1
X_12706_ _05173_ _05180_ VGND VGND VPWR VPWR _05182_ sky130_fd_sc_hd__and2_1
XFILLER_0_127_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10898_ _03134_ _03193_ VGND VGND VPWR VPWR _03194_ sky130_fd_sc_hd__nor2_1
X_13686_ _02427_ _02426_ _02735_ _02731_ VGND VGND VPWR VPWR _06242_ sky130_fd_sc_hd__and4_1
XFILLER_0_26_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07103__A _00486_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09021__C _00142_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12637_ _05105_ _05040_ VGND VGND VPWR VPWR _05106_ sky130_fd_sc_hd__nand2_1
XFILLER_0_143_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12568_ _05002_ _04996_ VGND VGND VPWR VPWR _05030_ sky130_fd_sc_hd__and2b_1
XFILLER_0_25_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11519_ _03868_ _03870_ VGND VGND VPWR VPWR _03876_ sky130_fd_sc_hd__nand2_2
XFILLER_0_123_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13478__C _01062_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12499_ _04947_ _04951_ _04953_ VGND VGND VPWR VPWR _04954_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_111_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14169_ _06743_ _06748_ _06767_ VGND VGND VPWR VPWR _06769_ sky130_fd_sc_hd__a21o_1
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10554__B1 _02723_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08730_ _00293_ VGND VGND VPWR VPWR _00819_ sky130_fd_sc_hd__clkbuf_4
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10857__A1 _05588_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09711__A2 _01508_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08661_ _00159_ _00742_ VGND VGND VPWR VPWR _00743_ sky130_fd_sc_hd__nand2_1
XANTENNA__10857__B2 _02304_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11445__D _03679_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07612_ _05967_ _05988_ _06054_ VGND VGND VPWR VPWR _06065_ sky130_fd_sc_hd__a21oi_2
X_08592_ _00469_ _00492_ _00490_ VGND VGND VPWR VPWR _00668_ sky130_fd_sc_hd__a21o_1
XFILLER_0_89_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07543_ _04807_ _04730_ VGND VGND VPWR VPWR _05324_ sky130_fd_sc_hd__or2b_1
XFILLER_0_88_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13271__A2 _05776_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07474_ _04411_ _04477_ _04554_ VGND VGND VPWR VPWR _04565_ sky130_fd_sc_hd__and3_1
XANTENNA__11461__C _01953_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08109__A _06417_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09213_ _01345_ _01346_ VGND VGND VPWR VPWR _01347_ sky130_fd_sc_hd__nor2_1
XFILLER_0_57_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11180__D _03503_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_146_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_168 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09144_ _01207_ _01214_ VGND VGND VPWR VPWR _01271_ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_138 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09075_ _01194_ _01195_ _01996_ net11 VGND VGND VPWR VPWR _01196_ sky130_fd_sc_hd__and4bb_1
XANTENNA__10374__A _06819_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11990__C1 _01958_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08026_ _00057_ _00068_ VGND VGND VPWR VPWR _00070_ sky130_fd_sc_hd__or2_1
XFILLER_0_114_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07386__C _03499_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07683__A net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09977_ _02183_ VGND VGND VPWR VPWR _02184_ sky130_fd_sc_hd__inv_2
XANTENNA__07961__A1 _02259_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07961__B2 _02171_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08928_ _00853_ _00856_ _01035_ VGND VGND VPWR VPWR _01036_ sky130_fd_sc_hd__a21oi_2
XANTENNA__10848__A1 _00541_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10848__B2 _05742_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08859_ _03587_ net47 _00959_ _03576_ VGND VGND VPWR VPWR _00960_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11870_ _06885_ _01780_ _04261_ VGND VGND VPWR VPWR _04262_ sky130_fd_sc_hd__and3_1
XFILLER_0_86_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10821_ _00891_ net56 net57 _00989_ VGND VGND VPWR VPWR _03109_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13540_ _06079_ _06080_ VGND VGND VPWR VPWR _06081_ sky130_fd_sc_hd__nor2_1
X_10752_ _02975_ _03032_ VGND VGND VPWR VPWR _03033_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_109_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12470__B1 _01289_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_375 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13471_ _05993_ _05989_ _06004_ VGND VGND VPWR VPWR _06005_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_82_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10683_ _02943_ _02944_ _02942_ VGND VGND VPWR VPWR _02957_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_125_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12422_ _04860_ _04868_ VGND VGND VPWR VPWR _04869_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12353_ _00742_ _00605_ _04791_ _04792_ VGND VGND VPWR VPWR _04793_ sky130_fd_sc_hd__a31o_1
XANTENNA__08441__A2 _00158_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09495__D net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11304_ _03638_ _03639_ VGND VGND VPWR VPWR _03640_ sky130_fd_sc_hd__and2_1
X_12284_ _04714_ _01182_ _04716_ VGND VGND VPWR VPWR _04717_ sky130_fd_sc_hd__a21o_1
XFILLER_0_10_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14023_ _05851_ _05421_ _05958_ VGND VGND VPWR VPWR _06612_ sky130_fd_sc_hd__o21a_1
XFILLER_0_120_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11235_ _03015_ _01062_ _01415_ _00410_ VGND VGND VPWR VPWR _03564_ sky130_fd_sc_hd__a22oi_1
X_11166_ _03458_ _03467_ VGND VGND VPWR VPWR _03489_ sky130_fd_sc_hd__nand2_1
X_10117_ _06937_ _02188_ VGND VGND VPWR VPWR _02337_ sky130_fd_sc_hd__nand2_1
X_11097_ _03409_ _03410_ VGND VGND VPWR VPWR _03413_ sky130_fd_sc_hd__and2_1
XANTENNA__12004__A _00257_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10048_ _02260_ _02261_ VGND VGND VPWR VPWR _02262_ sky130_fd_sc_hd__nor2_1
XFILLER_0_117_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13807_ _02190_ _03699_ _06367_ VGND VGND VPWR VPWR _06375_ sky130_fd_sc_hd__and3_1
XANTENNA__09457__A1 _06820_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09457__B2 net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11999_ _03990_ _03992_ VGND VGND VPWR VPWR _04404_ sky130_fd_sc_hd__nor2_2
XFILLER_0_133_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13738_ _05861_ _05866_ _06298_ VGND VGND VPWR VPWR _06299_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_128_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13669_ _06162_ _06222_ VGND VGND VPWR VPWR _06223_ sky130_fd_sc_hd__and2_1
XFILLER_0_45_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_414 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07190_ _01328_ _01427_ VGND VGND VPWR VPWR _01448_ sky130_fd_sc_hd__xor2_2
XFILLER_0_54_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09983__A _02189_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09900_ _01605_ _01786_ _01993_ _01991_ VGND VGND VPWR VPWR _02099_ sky130_fd_sc_hd__a31o_1
XFILLER_0_1_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09831_ _01771_ _02023_ VGND VGND VPWR VPWR _02024_ sky130_fd_sc_hd__xor2_1
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12315__A1_N _00608_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09762_ _01946_ _01945_ VGND VGND VPWR VPWR _01948_ sky130_fd_sc_hd__and2_2
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08713_ _00789_ _00799_ VGND VGND VPWR VPWR _00800_ sky130_fd_sc_hd__xnor2_1
X_09693_ _05192_ _00373_ _01701_ _01699_ VGND VGND VPWR VPWR _01872_ sky130_fd_sc_hd__a31o_1
XANTENNA__12849__A _01585_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xrebuffer11 _01985_ VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__clkbuf_2
XTAP_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08644_ _00721_ _00724_ VGND VGND VPWR VPWR _00725_ sky130_fd_sc_hd__and2_4
Xrebuffer22 _01164_ VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__clkbuf_1
Xrebuffer33 _02083_ VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08575_ _00642_ _00647_ VGND VGND VPWR VPWR _00649_ sky130_fd_sc_hd__and2_1
XTAP_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07526_ _00901_ _04378_ _05093_ _05126_ VGND VGND VPWR VPWR _05137_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_77_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07457_ _04367_ VGND VGND VPWR VPWR _04378_ sky130_fd_sc_hd__buf_4
XFILLER_0_147_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_356 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07388_ _03488_ _03609_ VGND VGND VPWR VPWR _03620_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10816__B _02731_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09127_ _02138_ _01182_ _01252_ _00344_ VGND VGND VPWR VPWR _01253_ sky130_fd_sc_hd__a22o_1
XANTENNA__12755__A1 _01180_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09058_ _01177_ VGND VGND VPWR VPWR _01178_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_142_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08009_ _00047_ _00052_ VGND VGND VPWR VPWR _00053_ sky130_fd_sc_hd__nor2_1
XANTENNA__08005__C _04367_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_686 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10832__A _01339_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11020_ _02558_ _03327_ VGND VGND VPWR VPWR _03328_ sky130_fd_sc_hd__nor2_1
XANTENNA__11191__B1 _01156_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12971_ _05430_ _05448_ VGND VGND VPWR VPWR _05473_ sky130_fd_sc_hd__xor2_2
XANTENNA__12759__A _00457_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11922_ _04212_ _04317_ _04316_ VGND VGND VPWR VPWR _04319_ sky130_fd_sc_hd__o21a_1
XFILLER_0_87_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11382__B _02249_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11853_ _04237_ _04241_ _04242_ VGND VGND VPWR VPWR _04243_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_86_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10279__A _01339_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10804_ _03085_ _03088_ VGND VGND VPWR VPWR _03090_ sky130_fd_sc_hd__or2_1
X_11784_ _04165_ _02657_ _04166_ VGND VGND VPWR VPWR _04167_ sky130_fd_sc_hd__and3_1
XFILLER_0_95_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13523_ _06036_ _06037_ _06060_ _06061_ VGND VGND VPWR VPWR _06062_ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10735_ _03008_ _03010_ _03013_ VGND VGND VPWR VPWR _03014_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_103_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13454_ _05985_ _02766_ VGND VGND VPWR VPWR _05986_ sky130_fd_sc_hd__nand2_1
X_10666_ _00819_ _00818_ _02856_ _02858_ VGND VGND VPWR VPWR _02939_ sky130_fd_sc_hd__and4_1
XFILLER_0_125_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12746__A1 _00378_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12405_ _04848_ _04849_ VGND VGND VPWR VPWR _04850_ sky130_fd_sc_hd__xnor2_1
X_13385_ _05899_ _05378_ _05909_ VGND VGND VPWR VPWR _05911_ sky130_fd_sc_hd__a21oi_1
X_10597_ _02859_ _02860_ _02854_ VGND VGND VPWR VPWR _02863_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_88_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09611__A1 _02335_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput109 net109 VGND VGND VPWR VPWR prod[4] sky130_fd_sc_hd__clkbuf_4
X_12336_ _04736_ _04773_ VGND VGND VPWR VPWR _04775_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_23_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12267_ _04661_ _04698_ VGND VGND VPWR VPWR _04699_ sky130_fd_sc_hd__xor2_2
XFILLER_0_120_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14006_ _06588_ _06589_ _06591_ VGND VGND VPWR VPWR _06594_ sky130_fd_sc_hd__and3_1
X_11218_ _03537_ _03544_ _03538_ VGND VGND VPWR VPWR _03546_ sky130_fd_sc_hd__or3_1
XANTENNA_output72_A net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09308__A _00844_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12198_ _04621_ _04612_ _04622_ VGND VGND VPWR VPWR _04623_ sky130_fd_sc_hd__o21a_1
Xoutput80 net80 VGND VGND VPWR VPWR prod[23] sky130_fd_sc_hd__clkbuf_4
Xoutput91 net91 VGND VGND VPWR VPWR prod[33] sky130_fd_sc_hd__clkbuf_4
X_11149_ _03042_ _03469_ VGND VGND VPWR VPWR _03470_ sky130_fd_sc_hd__nor2_2
XFILLER_0_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09127__B1 _01252_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12388__B _00779_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08360_ _00413_ VGND VGND VPWR VPWR _00414_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_58_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07311_ _02642_ _02653_ _02751_ VGND VGND VPWR VPWR _02773_ sky130_fd_sc_hd__nand3_2
XFILLER_0_46_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11788__A2 net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09697__B _04026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08291_ _00335_ _00338_ VGND VGND VPWR VPWR _00339_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07242_ _02007_ VGND VGND VPWR VPWR _02018_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14108__B _02743_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07173_ _01230_ _00672_ _01241_ _01251_ VGND VGND VPWR VPWR _01262_ sky130_fd_sc_hd__a31o_1
XFILLER_0_143_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09218__A _01311_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07916__A1 _01996_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09814_ _01610_ _01612_ _01803_ _02004_ VGND VGND VPWR VPWR _02005_ sky130_fd_sc_hd__a31o_4
X_09745_ _01918_ _01920_ _01927_ VGND VGND VPWR VPWR _01929_ sky130_fd_sc_hd__or3_1
XFILLER_0_94_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09676_ _01735_ _01852_ VGND VGND VPWR VPWR _01854_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07144__A2 net61 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08341__A1 _02138_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08341__B2 _00344_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08627_ _00666_ _00706_ VGND VGND VPWR VPWR _00707_ sky130_fd_sc_hd__xnor2_2
XTAP_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08558_ _00629_ _00630_ VGND VGND VPWR VPWR _00631_ sky130_fd_sc_hd__or2_1
XFILLER_0_77_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07509_ _00333_ _04917_ _04939_ _02138_ VGND VGND VPWR VPWR _04950_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08489_ _00181_ _00555_ _00346_ VGND VGND VPWR VPWR _00556_ sky130_fd_sc_hd__a21o_1
XFILLER_0_9_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10520_ _02772_ _02771_ VGND VGND VPWR VPWR _02778_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_64_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10451_ _02701_ _02702_ VGND VGND VPWR VPWR _02703_ sky130_fd_sc_hd__nand2_4
XFILLER_0_122_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08016__B _04510_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12837__A1_N _02728_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13170_ _05683_ _05689_ VGND VGND VPWR VPWR _05692_ sky130_fd_sc_hd__and2_1
X_10382_ _02623_ _02626_ VGND VGND VPWR VPWR _02627_ sky130_fd_sc_hd__nand2_1
X_12121_ _03956_ _04001_ VGND VGND VPWR VPWR _04538_ sky130_fd_sc_hd__and2_1
XFILLER_0_130_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12052_ _04244_ _04247_ _04249_ VGND VGND VPWR VPWR _04462_ sky130_fd_sc_hd__and3_1
X_11003_ _05192_ _04598_ _01368_ _00959_ VGND VGND VPWR VPWR _03309_ sky130_fd_sc_hd__and4_1
XANTENNA__07383__A2 _03554_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08580__A1 _00399_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08580__B2 _03015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12489__A _01517_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08686__B _04048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12954_ _05030_ _05003_ VGND VGND VPWR VPWR _05454_ sky130_fd_sc_hd__or2b_2
X_11905_ _04294_ _04297_ _04298_ _04296_ VGND VGND VPWR VPWR _04300_ sky130_fd_sc_hd__o22a_1
XANTENNA_output110_A net110 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12885_ _05243_ _05376_ VGND VGND VPWR VPWR _05378_ sky130_fd_sc_hd__nand2_1
XFILLER_0_114_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09798__A _03059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11836_ _04171_ _04192_ VGND VGND VPWR VPWR _04225_ sky130_fd_sc_hd__or2_1
XTAP_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08096__B1 _04928_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10737__A _00399_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11767_ _03070_ _02335_ _01954_ _02135_ VGND VGND VPWR VPWR _04149_ sky130_fd_sc_hd__and4_1
X_13506_ _06025_ _06028_ _06042_ VGND VGND VPWR VPWR _06044_ sky130_fd_sc_hd__a21oi_1
X_10718_ _02921_ _02923_ VGND VGND VPWR VPWR _02996_ sky130_fd_sc_hd__or2_1
XFILLER_0_70_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11698_ _04069_ _04071_ _04063_ _04065_ VGND VGND VPWR VPWR _04073_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_125_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__07111__A _00563_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12374__D _00607_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13437_ _05960_ _05968_ VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__xor2_4
XANTENNA__14184__A3 _06778_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xrebuffer2 _06932_ VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__buf_1
XFILLER_0_3_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10649_ _02796_ _02919_ VGND VGND VPWR VPWR _02920_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_24_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13368_ _05292_ _05353_ _05354_ _02765_ _02008_ VGND VGND VPWR VPWR _05893_ sky130_fd_sc_hd__a32o_1
X_12319_ _04753_ _04755_ VGND VGND VPWR VPWR _04756_ sky130_fd_sc_hd__and2b_1
XANTENNA__10472__A _02724_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13299_ _05694_ _05821_ VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__xnor2_4
XANTENNA__09038__A _00526_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07860_ _05401_ _06988_ VGND VGND VPWR VPWR _06989_ sky130_fd_sc_hd__nor2_1
X_07791_ _06916_ _06919_ VGND VGND VPWR VPWR _06920_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08596__B _06483_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09530_ _01539_ _01693_ VGND VGND VPWR VPWR _01694_ sky130_fd_sc_hd__and2_1
XFILLER_0_64_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07931__D net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09461_ _01617_ _03894_ _00475_ _01615_ VGND VGND VPWR VPWR _01619_ sky130_fd_sc_hd__and4b_1
XANTENNA__11453__D _03681_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08412_ _02149_ _00112_ _00268_ _05588_ VGND VGND VPWR VPWR _00471_ sky130_fd_sc_hd__a22o_1
X_09392_ _01064_ _01105_ _01406_ _01542_ VGND VGND VPWR VPWR _01543_ sky130_fd_sc_hd__a31o_1
XANTENNA__10681__A2 _01411_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08343_ _00384_ _00386_ _00395_ VGND VGND VPWR VPWR _00396_ sky130_fd_sc_hd__o21a_1
XFILLER_0_129_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13023__A _05509_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08274_ _00166_ _00169_ VGND VGND VPWR VPWR _00320_ sky130_fd_sc_hd__or2b_1
XFILLER_0_104_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08117__A _00157_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_116_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_570 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07225_ _01569_ _01810_ _01821_ VGND VGND VPWR VPWR _01832_ sky130_fd_sc_hd__o21bai_4
XFILLER_0_6_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_288 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07156_ _00869_ VGND VGND VPWR VPWR _01076_ sky130_fd_sc_hd__buf_4
XANTENNA__11933__A2 _00574_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07675__B _00989_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07087_ _00311_ VGND VGND VPWR VPWR _00322_ sky130_fd_sc_hd__buf_4
XFILLER_0_140_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07691__A net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07989_ _00019_ _00031_ VGND VGND VPWR VPWR _00033_ sky130_fd_sc_hd__or2_1
X_09728_ _01906_ _01909_ VGND VGND VPWR VPWR _01911_ sky130_fd_sc_hd__and2_1
XFILLER_0_69_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09659_ _01833_ _01834_ _01631_ VGND VGND VPWR VPWR _01836_ sky130_fd_sc_hd__a21o_1
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12670_ _04910_ _05035_ _04896_ VGND VGND VPWR VPWR _05142_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_139_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09411__A net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11621_ _00544_ _01182_ _03986_ VGND VGND VPWR VPWR _03988_ sky130_fd_sc_hd__and3_1
XFILLER_0_108_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11552_ _03904_ _03911_ VGND VGND VPWR VPWR _03912_ sky130_fd_sc_hd__or2b_1
XFILLER_0_92_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10276__B net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10503_ _02758_ VGND VGND VPWR VPWR _02759_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_108_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11483_ _03834_ _03835_ VGND VGND VPWR VPWR _03836_ sky130_fd_sc_hd__or2b_1
XFILLER_0_80_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13222_ _05628_ _05630_ _05748_ _05646_ VGND VGND VPWR VPWR _05749_ sky130_fd_sc_hd__a22o_1
X_10434_ _02447_ _02457_ VGND VGND VPWR VPWR _02684_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10365_ _02604_ _02607_ VGND VGND VPWR VPWR _02608_ sky130_fd_sc_hd__nand2_1
X_13153_ _05211_ _05672_ VGND VGND VPWR VPWR _05673_ sky130_fd_sc_hd__nand2_2
XFILLER_0_103_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12104_ _04492_ _04517_ _04518_ VGND VGND VPWR VPWR _04519_ sky130_fd_sc_hd__a21o_2
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13084_ _05506_ _05596_ _05505_ VGND VGND VPWR VPWR _05597_ sky130_fd_sc_hd__a21oi_2
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10296_ _02528_ _02531_ VGND VGND VPWR VPWR _02533_ sky130_fd_sc_hd__xor2_1
XANTENNA__11538__D _01564_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12035_ _04441_ _04374_ VGND VGND VPWR VPWR _04443_ sky130_fd_sc_hd__nand2_1
XFILLER_0_109_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11688__A1 _03510_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11688__B2 _00413_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08697__A _00782_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09305__B _01343_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11554__C _01177_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13986_ _06565_ _06570_ VGND VGND VPWR VPWR _06572_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07106__A _00519_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12937_ _04566_ _04582_ _04484_ VGND VGND VPWR VPWR _05436_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_88_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12868_ _05320_ _05321_ _05359_ VGND VGND VPWR VPWR _05360_ sky130_fd_sc_hd__a21o_1
XTAP_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11819_ _00157_ _03678_ _04205_ VGND VGND VPWR VPWR _04206_ sky130_fd_sc_hd__and3_1
XFILLER_0_145_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10467__A _02169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12799_ _05282_ _05283_ VGND VGND VPWR VPWR _05284_ sky130_fd_sc_hd__xnor2_1
XTAP_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11612__A1 _03554_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07479__C net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11612__B2 _00519_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13365__A1 _02765_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_64 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_792 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07595__A2 _05566_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08961_ _00963_ _00966_ _01070_ VGND VGND VPWR VPWR _01071_ sky130_fd_sc_hd__o21a_1
X_07912_ _02456_ _07040_ VGND VGND VPWR VPWR _07041_ sky130_fd_sc_hd__nand2_2
X_08892_ _03543_ _00144_ VGND VGND VPWR VPWR _00996_ sky130_fd_sc_hd__nand2_1
XANTENNA__12340__A2 _01368_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07843_ _06970_ _06971_ VGND VGND VPWR VPWR _06972_ sky130_fd_sc_hd__nand2_1
XANTENNA__08400__A _00457_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07774_ _01470_ net6 VGND VGND VPWR VPWR _06903_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09513_ _01672_ _01673_ _01670_ VGND VGND VPWR VPWR _01675_ sky130_fd_sc_hd__o21a_1
XFILLER_0_91_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09444_ _01586_ VGND VGND VPWR VPWR _01600_ sky130_fd_sc_hd__clkbuf_4
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09869__C _00755_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09375_ _01522_ _01523_ VGND VGND VPWR VPWR _01524_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10377__A _03521_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11911__D _03783_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12295__C _02190_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08326_ _04059_ VGND VGND VPWR VPWR _00378_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__10406__A2 _01564_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08257_ _00296_ _00301_ VGND VGND VPWR VPWR _00302_ sky130_fd_sc_hd__xnor2_2
XANTENNA__13688__A _02090_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07208_ _00891_ _00672_ VGND VGND VPWR VPWR _01645_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07686__A net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08188_ _00223_ _00216_ VGND VGND VPWR VPWR _00232_ sky130_fd_sc_hd__and2b_1
XANTENNA__10824__B _04268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_595 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07139_ _00880_ VGND VGND VPWR VPWR _00891_ sky130_fd_sc_hd__buf_6
XFILLER_0_113_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11001__A _02971_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10543__C _02724_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10150_ _02230_ _02371_ VGND VGND VPWR VPWR _02373_ sky130_fd_sc_hd__nor2_1
X_10081_ _02293_ VGND VGND VPWR VPWR _02297_ sky130_fd_sc_hd__inv_2
X_13840_ _06409_ _06410_ VGND VGND VPWR VPWR _06411_ sky130_fd_sc_hd__and2b_1
XANTENNA__11374__C _01957_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13771_ _06334_ VGND VGND VPWR VPWR _06335_ sky130_fd_sc_hd__inv_2
X_10983_ _03282_ _03285_ VGND VGND VPWR VPWR _03287_ sky130_fd_sc_hd__or2_1
XFILLER_0_139_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12722_ _00380_ _01182_ VGND VGND VPWR VPWR _05199_ sky130_fd_sc_hd__nand2_2
XFILLER_0_97_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08683__C _04015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12653_ _05122_ VGND VGND VPWR VPWR _05123_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11604_ _03958_ _03968_ VGND VGND VPWR VPWR _03969_ sky130_fd_sc_hd__and2_1
XFILLER_0_65_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12584_ _05045_ _05046_ VGND VGND VPWR VPWR _05047_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_26_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13598__A _01181_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11535_ _03778_ _03892_ VGND VGND VPWR VPWR _03893_ sky130_fd_sc_hd__and2_1
XANTENNA__09795__B _00138_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11466_ _03543_ _03681_ _03801_ _03802_ VGND VGND VPWR VPWR _03818_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_123_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13205_ _05722_ _05729_ VGND VGND VPWR VPWR _05730_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_111_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10417_ _02663_ _02665_ VGND VGND VPWR VPWR _02666_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11397_ _00112_ _01254_ _02119_ _00268_ VGND VGND VPWR VPWR _03742_ sky130_fd_sc_hd__a22o_1
X_14185_ _05960_ _06623_ _06643_ _06753_ VGND VGND VPWR VPWR _06784_ sky130_fd_sc_hd__or4_1
XFILLER_0_110_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13136_ _05652_ _05653_ VGND VGND VPWR VPWR _05655_ sky130_fd_sc_hd__nor2_1
X_10348_ _02382_ _02385_ _02588_ VGND VGND VPWR VPWR _02590_ sky130_fd_sc_hd__nand3_1
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_598 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11846__A _02456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10279_ _01339_ net53 VGND VGND VPWR VPWR _02514_ sky130_fd_sc_hd__nand2_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13067_ _02709_ _05578_ VGND VGND VPWR VPWR _05579_ sky130_fd_sc_hd__xnor2_4
X_12018_ _04423_ _04424_ VGND VGND VPWR VPWR _04425_ sky130_fd_sc_hd__nand2_1
XANTENNA__11565__B _02117_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08220__A _06472_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13969_ _06550_ _06552_ VGND VGND VPWR VPWR _06553_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07490_ net33 _04367_ VGND VGND VPWR VPWR _04741_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09160_ _01288_ VGND VGND VPWR VPWR _01289_ sky130_fd_sc_hd__buf_4
XANTENNA__12389__A2 _01586_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09201__D _00158_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08111_ _00055_ _00056_ _00053_ VGND VGND VPWR VPWR _00155_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_28_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09091_ _01212_ _01213_ VGND VGND VPWR VPWR _01214_ sky130_fd_sc_hd__nor2_1
XFILLER_0_114_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08042_ _00002_ _00085_ VGND VGND VPWR VPWR _00086_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_852 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09993_ _02198_ _02199_ VGND VGND VPWR VPWR _02201_ sky130_fd_sc_hd__and2_1
X_08944_ _01050_ _01052_ VGND VGND VPWR VPWR _01053_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_110_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12313__A2 _01601_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08875_ _00789_ _00799_ VGND VGND VPWR VPWR _00977_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07826_ _01076_ net37 VGND VGND VPWR VPWR _06955_ sky130_fd_sc_hd__nand2_1
X_07757_ _06848_ _06841_ VGND VGND VPWR VPWR _06886_ sky130_fd_sc_hd__or2b_1
XANTENNA__13813__A2 _03679_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07688_ _01120_ _03499_ _06813_ _06812_ VGND VGND VPWR VPWR _06817_ sky130_fd_sc_hd__a31o_1
XFILLER_0_66_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09427_ _01579_ _01581_ VGND VGND VPWR VPWR _01582_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09358_ _01368_ VGND VGND VPWR VPWR _01506_ sky130_fd_sc_hd__buf_2
XANTENNA__09245__A2 _00373_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08309_ _00240_ VGND VGND VPWR VPWR _00359_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09289_ _01429_ _01233_ _01430_ VGND VGND VPWR VPWR _01431_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_34_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12753__C _01248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11320_ _02917_ _03655_ _03657_ VGND VGND VPWR VPWR _03658_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_144_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_567 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11251_ _03580_ _03545_ _03581_ VGND VGND VPWR VPWR _03582_ sky130_fd_sc_hd__and3_1
XFILLER_0_120_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10202_ _02095_ _02429_ VGND VGND VPWR VPWR _02430_ sky130_fd_sc_hd__xor2_1
X_11182_ net138 _03505_ VGND VGND VPWR VPWR _03506_ sky130_fd_sc_hd__nor2_1
X_10133_ _02220_ _02221_ _02218_ VGND VGND VPWR VPWR _02354_ sky130_fd_sc_hd__a21o_1
XFILLER_0_101_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08508__A1 _02138_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08508__B2 _00333_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10064_ _02274_ _02278_ VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__xor2_2
XANTENNA__07582__C _00628_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10315__A1 _05192_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13823_ _05935_ _06391_ VGND VGND VPWR VPWR _06392_ sky130_fd_sc_hd__nor2_1
XANTENNA__12068__A1 _03554_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12068__B2 _00530_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13754_ _06299_ _06315_ VGND VGND VPWR VPWR _06316_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10966_ _03260_ _03267_ VGND VGND VPWR VPWR _03269_ sky130_fd_sc_hd__and2b_1
XFILLER_0_85_535 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12705_ _05177_ _05178_ _05179_ VGND VGND VPWR VPWR _05180_ sky130_fd_sc_hd__o21a_1
X_13685_ _06236_ _06239_ VGND VGND VPWR VPWR _06240_ sky130_fd_sc_hd__or2_1
X_10897_ _03133_ _03129_ _03131_ VGND VGND VPWR VPWR _03193_ sky130_fd_sc_hd__nor3_1
XFILLER_0_122_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12636_ _05102_ _05103_ VGND VGND VPWR VPWR _05105_ sky130_fd_sc_hd__xor2_1
XFILLER_0_26_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09021__D _04895_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12567_ _05018_ _05024_ _05026_ _05028_ VGND VGND VPWR VPWR _05029_ sky130_fd_sc_hd__o31ai_4
XFILLER_0_108_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11518_ _03868_ _03871_ _03874_ VGND VGND VPWR VPWR _03875_ sky130_fd_sc_hd__a21o_1
XFILLER_0_41_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08215__A _01383_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12498_ _04941_ _04952_ VGND VGND VPWR VPWR _04953_ sky130_fd_sc_hd__nor2_1
XFILLER_0_123_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11449_ _00262_ _03680_ _03798_ VGND VGND VPWR VPWR _03799_ sky130_fd_sc_hd__and3_1
XFILLER_0_111_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14168_ _06743_ _06748_ _06767_ VGND VGND VPWR VPWR _06768_ sky130_fd_sc_hd__and3_1
XFILLER_0_21_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10554__A1 _02993_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10554__B2 _00377_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11576__A _00262_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13119_ _04029_ _05635_ VGND VGND VPWR VPWR _05636_ sky130_fd_sc_hd__xnor2_4
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14099_ _06611_ _06693_ VGND VGND VPWR VPWR _06694_ sky130_fd_sc_hd__and2_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10857__A2 _01410_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08660_ _03773_ VGND VGND VPWR VPWR _00742_ sky130_fd_sc_hd__buf_4
X_07611_ _05999_ _06010_ _06043_ VGND VGND VPWR VPWR _06054_ sky130_fd_sc_hd__a21o_1
XFILLER_0_89_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08591_ _00493_ _00523_ VGND VGND VPWR VPWR _00667_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07542_ _00333_ _04939_ VGND VGND VPWR VPWR _05313_ sky130_fd_sc_hd__and2_2
XFILLER_0_72_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07473_ _04532_ _04543_ VGND VGND VPWR VPWR _04554_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11461__D _02134_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08109__B _00151_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09212_ _01149_ _01344_ VGND VGND VPWR VPWR _01346_ sky130_fd_sc_hd__and2_1
XFILLER_0_146_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09143_ _01206_ _01215_ VGND VGND VPWR VPWR _01270_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_810 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13031__A _05536_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09074_ _05445_ _00423_ net10 _05731_ VGND VGND VPWR VPWR _01195_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_112_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10793__A1 _06937_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10374__B _06821_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11990__B1 _00530_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08025_ _00057_ _00068_ VGND VGND VPWR VPWR _00069_ sky130_fd_sc_hd__nand2_1
XANTENNA__07386__D net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07683__B net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09976_ _02180_ _02181_ VGND VGND VPWR VPWR _02183_ sky130_fd_sc_hd__nand2_1
XANTENNA__07961__A2 _00004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08927_ _00673_ _00848_ _00852_ VGND VGND VPWR VPWR _01035_ sky130_fd_sc_hd__or3_1
X_08858_ net48 VGND VGND VPWR VPWR _00959_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07809_ _06626_ _06450_ _06937_ _06637_ VGND VGND VPWR VPWR _06938_ sky130_fd_sc_hd__and4_1
X_08789_ _00367_ _00554_ _00878_ _00879_ _00883_ VGND VGND VPWR VPWR _00884_ sky130_fd_sc_hd__o311a_4
XFILLER_0_67_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10820_ _03106_ _03107_ VGND VGND VPWR VPWR _03108_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_524 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07204__A _00420_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10751_ _02980_ _02983_ VGND VGND VPWR VPWR _03032_ sky130_fd_sc_hd__nor2_1
XANTENNA__12470__A1 _02008_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12470__B2 _04714_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13470_ _06002_ _06003_ VGND VGND VPWR VPWR _06004_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_387 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10682_ _02952_ _02955_ VGND VGND VPWR VPWR _02956_ sky130_fd_sc_hd__and2b_1
XFILLER_0_82_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12421_ _04866_ _04867_ VGND VGND VPWR VPWR _04868_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__08977__A1 _00541_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12483__C _00423_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__08977__B2 _00639_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12352_ _03696_ _03729_ _01506_ _01369_ VGND VGND VPWR VPWR _04792_ sky130_fd_sc_hd__and4_1
XFILLER_0_50_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11303_ _03629_ _03637_ VGND VGND VPWR VPWR _03639_ sky130_fd_sc_hd__or2_1
XFILLER_0_50_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12283_ _04715_ _04694_ VGND VGND VPWR VPWR _04716_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_132_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_660 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14022_ _05424_ _05960_ VGND VGND VPWR VPWR _06611_ sky130_fd_sc_hd__nor2_1
X_11234_ _03560_ _03561_ _03541_ VGND VGND VPWR VPWR _03563_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_30_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11396__A _00112_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11165_ _03484_ _03486_ VGND VGND VPWR VPWR _03487_ sky130_fd_sc_hd__and2_1
X_10116_ _02185_ _02197_ VGND VGND VPWR VPWR _02336_ sky130_fd_sc_hd__and2b_1
Xsplit3 _00869_ VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__buf_2
X_11096_ _03409_ _03410_ VGND VGND VPWR VPWR _03412_ sky130_fd_sc_hd__nor2_1
XANTENNA__12004__B _00670_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10047_ _02258_ _02245_ VGND VGND VPWR VPWR _02261_ sky130_fd_sc_hd__and2b_1
XFILLER_0_89_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13806_ _06366_ _06370_ _06372_ VGND VGND VPWR VPWR _06374_ sky130_fd_sc_hd__o21a_1
XFILLER_0_86_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11998_ _04401_ _04402_ VGND VGND VPWR VPWR _04403_ sky130_fd_sc_hd__nor2_4
XANTENNA__09457__A2 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13737_ _06293_ _06295_ VGND VGND VPWR VPWR _06298_ sky130_fd_sc_hd__xor2_1
X_10949_ _03108_ _03248_ _03249_ VGND VGND VPWR VPWR _03250_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_46_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13668_ _06152_ _06161_ _06160_ VGND VGND VPWR VPWR _06222_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_6_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12619_ _00415_ _00575_ _01060_ _01413_ VGND VGND VPWR VPWR _05086_ sky130_fd_sc_hd__and4_1
XFILLER_0_143_426 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13410__B1 _01956_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10475__A _02727_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13599_ _01061_ _03785_ _06144_ _06145_ _02856_ VGND VGND VPWR VPWR _06146_ sky130_fd_sc_hd__a32o_1
XFILLER_0_5_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13713__A1 _02427_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09917__B1 _01960_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13713__B2 _02726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09830_ _02021_ _02022_ VGND VGND VPWR VPWR _02023_ sky130_fd_sc_hd__and2b_1
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09761_ _01716_ _01717_ _01945_ _01946_ VGND VGND VPWR VPWR _01947_ sky130_fd_sc_hd__a211oi_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13477__B1 _03687_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08712_ _00797_ _00798_ VGND VGND VPWR VPWR _00799_ sky130_fd_sc_hd__or2_1
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09692_ _01703_ _01707_ VGND VGND VPWR VPWR _01871_ sky130_fd_sc_hd__nor2_1
XANTENNA__12849__B _01060_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xrebuffer12 _07060_ VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__clkbuf_1
X_08643_ _00565_ _00566_ _00569_ _00723_ VGND VGND VPWR VPWR _00724_ sky130_fd_sc_hd__o31ai_1
Xrebuffer23 net168 VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__clkbuf_1
Xrebuffer34 _04977_ VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__dlymetal6s4s_1
XFILLER_0_13_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08574_ _00642_ _00647_ VGND VGND VPWR VPWR _00648_ sky130_fd_sc_hd__nor2_1
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_332 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07525_ _05104_ VGND VGND VPWR VPWR _05126_ sky130_fd_sc_hd__inv_2
XFILLER_0_119_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07959__A _06765_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07456_ net2 VGND VGND VPWR VPWR _04367_ sky130_fd_sc_hd__buf_6
XFILLER_0_9_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07387_ _03565_ _03598_ VGND VGND VPWR VPWR _03609_ sky130_fd_sc_hd__or2_2
XFILLER_0_91_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09126_ _01250_ VGND VGND VPWR VPWR _01252_ sky130_fd_sc_hd__buf_4
XFILLER_0_115_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_610 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09057_ net17 VGND VGND VPWR VPWR _01177_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_142_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08008_ _00050_ _00051_ VGND VGND VPWR VPWR _00052_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10832__B net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09959_ _02154_ _02162_ VGND VGND VPWR VPWR _02164_ sky130_fd_sc_hd__nand2_1
X_12970_ _05453_ _05471_ VGND VGND VPWR VPWR _05472_ sky130_fd_sc_hd__xor2_4
XFILLER_0_99_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11921_ _04316_ _04212_ _04317_ VGND VGND VPWR VPWR _04318_ sky130_fd_sc_hd__nor3_1
XANTENNA__09414__A _04510_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11852_ _02663_ _04238_ _04240_ VGND VGND VPWR VPWR _04242_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10279__B net53 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10803_ _03085_ _03088_ VGND VGND VPWR VPWR _03089_ sky130_fd_sc_hd__nand2_1
X_11783_ _04151_ _04156_ VGND VGND VPWR VPWR _04166_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_55_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13522_ _06009_ _06018_ _03697_ _03699_ VGND VGND VPWR VPWR _06061_ sky130_fd_sc_hd__nand4_1
X_10734_ _02887_ _03012_ VGND VGND VPWR VPWR _03013_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13453_ _03783_ VGND VGND VPWR VPWR _05985_ sky130_fd_sc_hd__buf_2
XFILLER_0_36_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10665_ _02838_ _02936_ VGND VGND VPWR VPWR _02937_ sky130_fd_sc_hd__nor2_1
XFILLER_0_70_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12404_ _00374_ _01272_ VGND VGND VPWR VPWR _04849_ sky130_fd_sc_hd__nand2_1
XANTENNA__12746__A2 _03681_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_651 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13384_ _05899_ _05378_ _05909_ VGND VGND VPWR VPWR _05910_ sky130_fd_sc_hd__and3_1
XFILLER_0_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10596_ _02854_ _02859_ _02860_ VGND VGND VPWR VPWR _02862_ sky130_fd_sc_hd__and3_1
XANTENNA__09611__A2 _01780_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12335_ _04744_ _04746_ _04772_ VGND VGND VPWR VPWR _04773_ sky130_fd_sc_hd__a21o_1
XFILLER_0_133_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12266_ _04673_ _04696_ _04671_ VGND VGND VPWR VPWR _04698_ sky130_fd_sc_hd__a21o_1
X_14005_ _06590_ _06591_ VGND VGND VPWR VPWR _06592_ sky130_fd_sc_hd__nor2_1
XANTENNA__08178__A2 _00219_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11217_ _03537_ _03538_ _03544_ VGND VGND VPWR VPWR _03545_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_120_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09308__B _00819_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput70 net70 VGND VGND VPWR VPWR prod[14] sky130_fd_sc_hd__clkbuf_4
X_12197_ _03453_ _03468_ _03492_ VGND VGND VPWR VPWR _04622_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_120_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput81 net81 VGND VGND VPWR VPWR prod[24] sky130_fd_sc_hd__clkbuf_4
Xoutput92 net92 VGND VGND VPWR VPWR prod[34] sky130_fd_sc_hd__clkbuf_4
XANTENNA__07109__A net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11148_ _03038_ _03040_ _03031_ VGND VGND VPWR VPWR _03469_ sky130_fd_sc_hd__o21a_1
XANTENNA__09127__A1 _02138_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09127__B2 _00344_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11079_ _03361_ _03392_ VGND VGND VPWR VPWR _03393_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09324__A _00844_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12388__C _01586_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10189__B _00734_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07310_ _02642_ _02653_ _02751_ VGND VGND VPWR VPWR _02762_ sky130_fd_sc_hd__a21oi_1
X_08290_ _00336_ _00337_ VGND VGND VPWR VPWR _00338_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07241_ _01996_ VGND VGND VPWR VPWR _02007_ sky130_fd_sc_hd__buf_4
XFILLER_0_144_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07172_ net176 net149 _00705_ _00573_ VGND VGND VPWR VPWR _01251_ sky130_fd_sc_hd__and4_1
XFILLER_0_54_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08403__A _00453_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13698__B1 _02730_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09218__B _01352_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07916__A2 _04378_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09813_ _01804_ _01801_ _01802_ VGND VGND VPWR VPWR _02004_ sky130_fd_sc_hd__o21ai_1
X_09744_ _01918_ _01920_ _01927_ VGND VGND VPWR VPWR _01928_ sky130_fd_sc_hd__o21a_1
X_09675_ _01850_ _01851_ VGND VGND VPWR VPWR _01852_ sky130_fd_sc_hd__nor2_1
XTAP_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08341__A2 _00391_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08626_ _00667_ _00704_ VGND VGND VPWR VPWR _00706_ sky130_fd_sc_hd__xor2_1
XTAP_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08557_ _00599_ _00600_ _00627_ VGND VGND VPWR VPWR _00630_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_37_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07689__A net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07508_ _04928_ VGND VGND VPWR VPWR _04939_ sky130_fd_sc_hd__buf_4
XFILLER_0_147_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08488_ _00252_ _00253_ _00343_ VGND VGND VPWR VPWR _00555_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_91_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10987__A1 _00310_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_595 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07439_ net42 VGND VGND VPWR VPWR _04180_ sky130_fd_sc_hd__buf_2
XFILLER_0_80_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10450_ _02699_ _02700_ VGND VGND VPWR VPWR _02702_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_755 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09109_ _01176_ _01233_ VGND VGND VPWR VPWR _01234_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_60_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08016__C net6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_115_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10381_ _02624_ _02625_ VGND VGND VPWR VPWR _02626_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_32_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12120_ _04531_ _04536_ VGND VGND VPWR VPWR _04537_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12051_ _04459_ _04460_ VGND VGND VPWR VPWR _04461_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11002_ _05181_ _00604_ _03306_ _03307_ VGND VGND VPWR VPWR _03308_ sky130_fd_sc_hd__a31oi_2
XANTENNA__08580__A2 _00654_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13592__C _01414_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12489__B _00916_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12953_ _05449_ _05451_ _05452_ VGND VGND VPWR VPWR _05453_ sky130_fd_sc_hd__a21o_2
XFILLER_0_87_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11904_ _04294_ _04296_ _04297_ _04298_ VGND VGND VPWR VPWR _04299_ sky130_fd_sc_hd__nor4_1
XTAP_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12884_ _05243_ _05376_ VGND VGND VPWR VPWR _05377_ sky130_fd_sc_hd__or2_1
XTAP_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11835_ _04219_ _04222_ VGND VGND VPWR VPWR _04223_ sky130_fd_sc_hd__nor2_1
XFILLER_0_114_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output103_A net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09798__B _01585_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08096__A1 _02018_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08096__B2 _05478_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_110 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11766_ _04145_ _04146_ VGND VGND VPWR VPWR _04148_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_56_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10737__B _03015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13505_ _06040_ _06041_ VGND VGND VPWR VPWR _06042_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10717_ _02991_ _02994_ VGND VGND VPWR VPWR _02995_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11697_ _04063_ _04065_ _04069_ _04071_ VGND VGND VPWR VPWR _04072_ sky130_fd_sc_hd__o211a_1
XFILLER_0_126_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07111__B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13436_ _05833_ _05962_ _05966_ VGND VGND VPWR VPWR _05968_ sky130_fd_sc_hd__a21oi_4
X_10648_ _02917_ _02918_ VGND VGND VPWR VPWR _02919_ sky130_fd_sc_hd__nor2_2
XFILLER_0_141_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrebuffer3 _01810_ VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_63_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09596__A1 _00475_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13367_ _05292_ _05354_ _05353_ VGND VGND VPWR VPWR _05892_ sky130_fd_sc_hd__a21o_1
XFILLER_0_106_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10579_ _00143_ _04906_ _02306_ _02305_ VGND VGND VPWR VPWR _02843_ sky130_fd_sc_hd__and4_1
XFILLER_0_23_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12318_ _04750_ _04754_ VGND VGND VPWR VPWR _04755_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13298_ _05777_ _05794_ _05815_ _05816_ _05820_ VGND VGND VPWR VPWR _05821_ sky130_fd_sc_hd__o311a_4
XANTENNA__09348__A1 _00612_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12249_ _04663_ _04662_ VGND VGND VPWR VPWR _04679_ sky130_fd_sc_hd__or2b_1
XFILLER_0_139_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07790_ _06917_ _06918_ VGND VGND VPWR VPWR _06919_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08596__C _00113_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08859__B1 _00959_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09460_ _00475_ _03894_ _01616_ _01617_ VGND VGND VPWR VPWR _01618_ sky130_fd_sc_hd__o2bb2a_1
X_08411_ _06494_ _07004_ _00274_ _00277_ VGND VGND VPWR VPWR _00470_ sky130_fd_sc_hd__a31o_1
XFILLER_0_59_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_652 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09391_ _01403_ _01404_ VGND VGND VPWR VPWR _01542_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08342_ _03751_ _00394_ VGND VGND VPWR VPWR _00395_ sky130_fd_sc_hd__nor2_2
XFILLER_0_47_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_584 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08273_ _00303_ _00318_ VGND VGND VPWR VPWR _00319_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08117__B _00158_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07224_ _01536_ _01558_ VGND VGND VPWR VPWR _01821_ sky130_fd_sc_hd__and2b_1
XFILLER_0_73_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13958__B _06540_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07155_ _01033_ _01055_ VGND VGND VPWR VPWR _01065_ sky130_fd_sc_hd__and2b_1
XFILLER_0_70_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__14135__A _02743_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__12591__B1 _02857_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07086_ _00300_ VGND VGND VPWR VPWR _00311_ sky130_fd_sc_hd__buf_4
XANTENNA__07675__C _06733_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12343__B1 _01369_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07988_ _00019_ _00031_ VGND VGND VPWR VPWR _00032_ sky130_fd_sc_hd__nand2_1
X_09727_ _01906_ _01909_ VGND VGND VPWR VPWR _01910_ sky130_fd_sc_hd__nor2_1
XFILLER_0_69_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09511__A1 _06494_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10657__B1 _02722_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09658_ _01631_ _01833_ _01834_ VGND VGND VPWR VPWR _01835_ sky130_fd_sc_hd__nand3_1
XFILLER_0_69_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08609_ _00496_ _00522_ _00520_ VGND VGND VPWR VPWR _00687_ sky130_fd_sc_hd__a21o_1
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09589_ _01718_ _01754_ _01758_ VGND VGND VPWR VPWR _01759_ sky130_fd_sc_hd__and3_1
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_836 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11620_ _00544_ _01182_ _03986_ VGND VGND VPWR VPWR _03987_ sky130_fd_sc_hd__a21o_1
XFILLER_0_37_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11551_ _03909_ _03910_ VGND VGND VPWR VPWR _03911_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10502_ _01934_ VGND VGND VPWR VPWR _02758_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_135_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11482_ _03808_ _03810_ VGND VGND VPWR VPWR _03835_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_80_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13221_ _05644_ VGND VGND VPWR VPWR _05748_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10433_ _02666_ _02682_ VGND VGND VPWR VPWR _02683_ sky130_fd_sc_hd__xor2_1
XFILLER_0_116_790 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13152_ _05182_ VGND VGND VPWR VPWR _05672_ sky130_fd_sc_hd__inv_2
X_10364_ _02605_ _02606_ VGND VGND VPWR VPWR _02607_ sky130_fd_sc_hd__xnor2_1
X_12103_ _04515_ _04516_ VGND VGND VPWR VPWR _04518_ sky130_fd_sc_hd__nor2_1
XFILLER_0_103_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13083_ _05519_ _05523_ VGND VGND VPWR VPWR _05596_ sky130_fd_sc_hd__or2_1
X_10295_ _02529_ _02530_ VGND VGND VPWR VPWR _02531_ sky130_fd_sc_hd__xnor2_1
X_12034_ _04441_ _04374_ VGND VGND VPWR VPWR _04442_ sky130_fd_sc_hd__or2_1
XANTENNA__11688__A2 _00734_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13985_ _06568_ _06569_ VGND VGND VPWR VPWR _06570_ sky130_fd_sc_hd__nor2_1
X_12936_ _05433_ VGND VGND VPWR VPWR _05435_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12867_ _05356_ _05358_ VGND VGND VPWR VPWR _05359_ sky130_fd_sc_hd__xnor2_1
XTAP_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11818_ _00159_ _03682_ VGND VGND VPWR VPWR _04205_ sky130_fd_sc_hd__nand2_1
XANTENNA__08218__A _06965_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12798_ _00916_ _01933_ VGND VGND VPWR VPWR _05283_ sky130_fd_sc_hd__nand2_1
XTAP_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07122__A net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07816__A1 net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11612__A2 _01956_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_508 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11749_ _04109_ _04112_ VGND VGND VPWR VPWR _04129_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_316 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13419_ _01183_ _01415_ _01252_ _01108_ VGND VGND VPWR VPWR _05949_ sky130_fd_sc_hd__a22o_1
XANTENNA__10483__A _02731_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_248 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08960_ _00964_ _00965_ VGND VGND VPWR VPWR _01070_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07911_ _04939_ VGND VGND VPWR VPWR _07040_ sky130_fd_sc_hd__buf_4
X_08891_ _00993_ _00994_ VGND VGND VPWR VPWR _00995_ sky130_fd_sc_hd__and2b_1
X_07842_ _06967_ _06968_ _06969_ _06963_ VGND VGND VPWR VPWR _06971_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_75_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07773_ _06900_ _06901_ VGND VGND VPWR VPWR _06902_ sky130_fd_sc_hd__and2b_1
XANTENNA__13018__B _05507_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09512_ _01670_ _01672_ _01673_ VGND VGND VPWR VPWR _01674_ sky130_fd_sc_hd__nor3_1
XFILLER_0_78_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09443_ _00416_ _01597_ _01598_ VGND VGND VPWR VPWR _01599_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_78_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09869__D _00741_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09374_ _01388_ _01391_ _01521_ VGND VGND VPWR VPWR _01523_ sky130_fd_sc_hd__nor3_1
XFILLER_0_136_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__10377__B _00734_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12295__D _02088_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08325_ _00375_ VGND VGND VPWR VPWR _00376_ sky130_fd_sc_hd__buf_4
XFILLER_0_145_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12873__A _00458_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__07967__A _00891_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08256_ _00061_ _00161_ _00297_ _00299_ VGND VGND VPWR VPWR _00301_ sky130_fd_sc_hd__a211o_1
XANTENNA__13688__B _02725_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07207_ _01514_ _01503_ VGND VGND VPWR VPWR _01635_ sky130_fd_sc_hd__and2b_1
XANTENNA__07686__B net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08187_ _02949_ _03631_ _00229_ _00230_ VGND VGND VPWR VPWR _00231_ sky130_fd_sc_hd__a31o_1
XFILLER_0_104_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07138_ _00869_ VGND VGND VPWR VPWR _00880_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_70_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11001__B _04378_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10543__D _02727_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10080_ _01443_ _01444_ _02294_ _02295_ _01486_ VGND VGND VPWR VPWR _02296_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_100_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__14069__B1 _02742_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11374__D _03690_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13770_ _06332_ _06333_ VGND VGND VPWR VPWR _06334_ sky130_fd_sc_hd__and2_1
X_10982_ _03282_ _03285_ VGND VGND VPWR VPWR _03286_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09422__A _06428_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12721_ _00391_ _01108_ _05197_ VGND VGND VPWR VPWR _05198_ sky130_fd_sc_hd__nand3_1
XFILLER_0_84_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09779__D net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12652_ _00390_ _02759_ _05121_ VGND VGND VPWR VPWR _05122_ sky130_fd_sc_hd__and3_1
XFILLER_0_37_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11603_ _03964_ _03966_ _03967_ VGND VGND VPWR VPWR _03968_ sky130_fd_sc_hd__o21a_1
XFILLER_0_38_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12583_ _00745_ _01412_ VGND VGND VPWR VPWR _05046_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11534_ _03776_ _03777_ VGND VGND VPWR VPWR _03892_ sky130_fd_sc_hd__or2_1
XANTENNA__13598__B _01413_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09795__C _00572_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_524 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11399__A _02120_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11465_ _03814_ _03815_ _03812_ VGND VGND VPWR VPWR _03816_ sky130_fd_sc_hd__o21ai_1
X_13204_ _05717_ _05718_ VGND VGND VPWR VPWR _05729_ sky130_fd_sc_hd__xnor2_1
X_10416_ _02646_ _02442_ _02647_ _02662_ VGND VGND VPWR VPWR _02665_ sky130_fd_sc_hd__o31ai_2
X_14184_ _06771_ _06776_ _06778_ _06781_ _06783_ VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__a311o_1
XFILLER_0_0_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11396_ _00112_ _00268_ _01254_ _02119_ VGND VGND VPWR VPWR _03741_ sky130_fd_sc_hd__and4_1
XFILLER_0_60_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13135_ _05634_ _05636_ VGND VGND VPWR VPWR _05653_ sky130_fd_sc_hd__xor2_2
X_10347_ _02382_ _02385_ _02588_ VGND VGND VPWR VPWR _02589_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11846__B _01955_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13066_ _05569_ _05576_ VGND VGND VPWR VPWR _05578_ sky130_fd_sc_hd__xnor2_4
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10278_ _01372_ net53 _02314_ _02172_ _02312_ VGND VGND VPWR VPWR _02513_ sky130_fd_sc_hd__a32o_1
X_12017_ _04421_ _04346_ VGND VGND VPWR VPWR _04424_ sky130_fd_sc_hd__nand2_1
XANTENNA__08220__B _06483_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07117__A _00639_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap1 _03504_ VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__clkbuf_1
XANTENNA__13283__A1 _05786_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13968_ _06475_ _06551_ VGND VGND VPWR VPWR _06552_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12919_ _05414_ _05415_ VGND VGND VPWR VPWR _05416_ sky130_fd_sc_hd__xnor2_2
X_13899_ _06470_ _06475_ VGND VGND VPWR VPWR _06476_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_622 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_400 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08110_ _00050_ _00153_ VGND VGND VPWR VPWR _00154_ sky130_fd_sc_hd__xor2_1
XFILLER_0_84_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09090_ _01744_ _01211_ _01209_ _01210_ VGND VGND VPWR VPWR _01213_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_142_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08041_ _00083_ _00084_ VGND VGND VPWR VPWR _00085_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12546__B1 _01400_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09992_ _02198_ _02199_ VGND VGND VPWR VPWR _02200_ sky130_fd_sc_hd__nor2_1
X_08943_ _01051_ VGND VGND VPWR VPWR _01052_ sky130_fd_sc_hd__inv_2
XANTENNA__09507__A _06472_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09714__A1 _06494_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08874_ _00957_ _00975_ VGND VGND VPWR VPWR _00976_ sky130_fd_sc_hd__xnor2_2
X_07825_ _06952_ _06953_ VGND VGND VPWR VPWR _06954_ sky130_fd_sc_hd__and2b_1
X_07756_ _06775_ VGND VGND VPWR VPWR _06885_ sky130_fd_sc_hd__buf_4
XANTENNA__13274__A1 _05784_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07687_ _06814_ _06815_ VGND VGND VPWR VPWR _06816_ sky130_fd_sc_hd__xnor2_1
Xsplit17 _00716_ VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__buf_6
X_09426_ _01574_ _01267_ _01578_ VGND VGND VPWR VPWR _01581_ sky130_fd_sc_hd__or3_1
XFILLER_0_94_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09357_ _01504_ VGND VGND VPWR VPWR _01505_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_35_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08308_ _00356_ _00357_ VGND VGND VPWR VPWR _00358_ sky130_fd_sc_hd__or2_1
XFILLER_0_90_731 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09288_ _01112_ _01174_ VGND VGND VPWR VPWR _01430_ sky130_fd_sc_hd__nor2_1
XFILLER_0_133_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08239_ _00267_ _00282_ VGND VGND VPWR VPWR _00283_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_50_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11250_ _03537_ _03544_ _03538_ _03547_ VGND VGND VPWR VPWR _03581_ sky130_fd_sc_hd__o31ai_2
XFILLER_0_105_579 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10201_ _06626_ _02426_ _02428_ VGND VGND VPWR VPWR _02429_ sky130_fd_sc_hd__and3_1
XANTENNA__09953__A1 _04268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09953__B2 _01372_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11181_ _03475_ _03480_ VGND VGND VPWR VPWR _03505_ sky130_fd_sc_hd__xor2_2
XANTENNA__10851__A _02664_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10132_ _02350_ _02352_ VGND VGND VPWR VPWR _02353_ sky130_fd_sc_hd__xor2_2
XANTENNA__08508__A2 _00415_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10063_ _01433_ _01437_ _01636_ _02275_ _02277_ VGND VGND VPWR VPWR _02278_ sky130_fd_sc_hd__a41o_2
XANTENNA__07582__D _05742_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10315__A2 net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13822_ _06389_ _06390_ VGND VGND VPWR VPWR _06391_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13265__A1 _05507_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12068__A2 _01183_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13753_ _05861_ _05866_ _06298_ VGND VGND VPWR VPWR _06315_ sky130_fd_sc_hd__or3_1
X_10965_ _03265_ _03266_ VGND VGND VPWR VPWR _03267_ sky130_fd_sc_hd__and2_1
X_12704_ _05174_ _05176_ VGND VGND VPWR VPWR _05179_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13684_ _06189_ _06235_ VGND VGND VPWR VPWR _06239_ sky130_fd_sc_hd__and2_1
X_10896_ _03176_ _03190_ VGND VGND VPWR VPWR _03192_ sky130_fd_sc_hd__xor2_1
XFILLER_0_85_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12635_ _00915_ _01933_ VGND VGND VPWR VPWR _05103_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_107 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12566_ _05017_ _05014_ VGND VGND VPWR VPWR _05028_ sky130_fd_sc_hd__or2b_1
XFILLER_0_31_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_135 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__07400__A _02127_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11517_ _03855_ _03873_ VGND VGND VPWR VPWR _03874_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13121__B _05620_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12497_ _04938_ _04940_ _04937_ VGND VGND VPWR VPWR _04952_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08215__B _01350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output95_A net95 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11448_ _00263_ _03683_ VGND VGND VPWR VPWR _03798_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10003__A1 _05181_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14167_ _06763_ _06766_ VGND VGND VPWR VPWR _06767_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11379_ _03711_ _03712_ _03721_ VGND VGND VPWR VPWR _03722_ sky130_fd_sc_hd__or3_1
XFILLER_0_21_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10554__A2 _02168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13118_ _05609_ _05615_ _05617_ _04031_ VGND VGND VPWR VPWR _05635_ sky130_fd_sc_hd__o31a_2
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09327__A _00145_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11576__B _03748_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08231__A _05566_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14098_ _06619_ _06632_ VGND VGND VPWR VPWR _06693_ sky130_fd_sc_hd__nor2_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13049_ _04971_ _05558_ VGND VGND VPWR VPWR _05559_ sky130_fd_sc_hd__nor2_4
XFILLER_0_147_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_820 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07610_ _05999_ _06010_ _06032_ VGND VGND VPWR VPWR _06043_ sky130_fd_sc_hd__o21a_1
X_08590_ _00664_ _00665_ VGND VGND VPWR VPWR _00666_ sky130_fd_sc_hd__or2_2
XFILLER_0_89_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09062__A _01181_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07541_ _04983_ _05291_ VGND VGND VPWR VPWR _05302_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07472_ _04499_ _04521_ _04488_ VGND VGND VPWR VPWR _04543_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09880__B1 _01288_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09211_ _01149_ _01344_ VGND VGND VPWR VPWR _01345_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07628__A1_N _02007_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09142_ _01267_ _01268_ VGND VGND VPWR VPWR _01269_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_658 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_822 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09073_ _05445_ _05731_ _03718_ net10 VGND VGND VPWR VPWR _01194_ sky130_fd_sc_hd__and4_1
XFILLER_0_72_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10793__A2 _02758_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10374__C _00730_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08024_ _00066_ _00067_ VGND VGND VPWR VPWR _00068_ sky130_fd_sc_hd__xor2_1
XFILLER_0_114_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11767__A _03070_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09975_ _02153_ _02179_ VGND VGND VPWR VPWR _02181_ sky130_fd_sc_hd__nand2_1
XANTENNA__07683__C net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08926_ _00857_ _00871_ VGND VGND VPWR VPWR _01034_ sky130_fd_sc_hd__and2_1
X_08857_ _00431_ _04169_ net47 net48 VGND VGND VPWR VPWR _00958_ sky130_fd_sc_hd__and4_1
XFILLER_0_99_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12598__A _03707_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07808_ _06472_ VGND VGND VPWR VPWR _06937_ sky130_fd_sc_hd__buf_4
X_08788_ _00711_ _00881_ _00882_ VGND VGND VPWR VPWR _00883_ sky130_fd_sc_hd__a21o_1
XFILLER_0_79_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07739_ _01284_ _06744_ VGND VGND VPWR VPWR _06868_ sky130_fd_sc_hd__nand2_1
XANTENNA__11007__A _00293_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__07204__B _00978_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10750_ _03029_ _03030_ VGND VGND VPWR VPWR _03031_ sky130_fd_sc_hd__or2_1
XFILLER_0_94_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12470__A2 _03414_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09409_ _01298_ _01299_ _01303_ VGND VGND VPWR VPWR _01562_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10681_ _00094_ _01411_ _02953_ _02954_ VGND VGND VPWR VPWR _02955_ sky130_fd_sc_hd__a31o_1
XFILLER_0_82_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_399 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12420_ _04850_ _04856_ VGND VGND VPWR VPWR _04867_ sky130_fd_sc_hd__xor2_1
XFILLER_0_35_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_800 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12483__D _03762_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12351_ _03729_ _01506_ _01369_ _03696_ VGND VGND VPWR VPWR _04791_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11302_ _03629_ _03637_ VGND VGND VPWR VPWR _03638_ sky130_fd_sc_hd__nand2_1
X_12282_ _04695_ _04687_ VGND VGND VPWR VPWR _04715_ sky130_fd_sc_hd__or2b_1
XFILLER_0_105_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14021_ _06238_ _06609_ VGND VGND VPWR VPWR _06610_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_132_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11233_ _03560_ _03541_ _03561_ VGND VGND VPWR VPWR _03562_ sky130_fd_sc_hd__and3_1
XANTENNA__09147__A _01361_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11164_ _03464_ _03485_ VGND VGND VPWR VPWR _03486_ sky130_fd_sc_hd__xnor2_4
XANTENNA__11396__B _00268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08051__A _00094_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10115_ _02180_ _02333_ VGND VGND VPWR VPWR _02334_ sky130_fd_sc_hd__xor2_2
X_11095_ _03391_ _03393_ VGND VGND VPWR VPWR _03410_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12004__C _02090_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07890__A _02719_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10046_ _02245_ _02258_ VGND VGND VPWR VPWR _02260_ sky130_fd_sc_hd__and2b_1
XFILLER_0_117_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_138 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13805_ _06365_ _06371_ VGND VGND VPWR VPWR _06372_ sky130_fd_sc_hd__nor2_1
X_11997_ _04398_ _04399_ _04328_ VGND VGND VPWR VPWR _04402_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_98_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__12997__B1 _05501_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10948_ _03064_ _03067_ _03104_ _03106_ _03065_ VGND VGND VPWR VPWR _03249_ sky130_fd_sc_hd__a311o_1
X_13736_ _06293_ _06295_ VGND VGND VPWR VPWR _06297_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09610__A _02280_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13667_ _01108_ _06075_ VGND VGND VPWR VPWR _06221_ sky130_fd_sc_hd__nand2_1
X_10879_ _03168_ _03171_ VGND VGND VPWR VPWR _03173_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12618_ _05041_ _05042_ _05084_ VGND VGND VPWR VPWR _05085_ sky130_fd_sc_hd__a21oi_1
X_13598_ _01181_ _01413_ _01250_ VGND VGND VPWR VPWR _06145_ sky130_fd_sc_hd__and3_1
XANTENNA__13410__B2 _04714_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__07130__A net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_143_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12549_ _05008_ net185 VGND VGND VPWR VPWR _05009_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09917__A1 _01361_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14219_ _06804_ VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__clkbuf_1
XANTENNA__13713__A2 _02758_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09917__B2 _00159_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09057__A net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09760_ _01713_ _01715_ VGND VGND VPWR VPWR _01946_ sky130_fd_sc_hd__nor2_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13477__B2 _01414_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08711_ _00790_ _00796_ VGND VGND VPWR VPWR _00798_ sky130_fd_sc_hd__nor2_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09691_ _05181_ _04059_ _01705_ VGND VGND VPWR VPWR _01870_ sky130_fd_sc_hd__and3_1
X_08642_ _00565_ _00722_ VGND VGND VPWR VPWR _00723_ sky130_fd_sc_hd__xnor2_1
Xrebuffer13 _07060_ VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__clkbuf_1
Xrebuffer24 _04697_ VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__clkbuf_1
XANTENNA__12211__A _00376_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xrebuffer35 _04596_ VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__buf_6
XFILLER_0_83_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08573_ _00643_ _00646_ VGND VGND VPWR VPWR _00647_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07524_ _05093_ _05104_ _00901_ _04378_ VGND VGND VPWR VPWR _05115_ sky130_fd_sc_hd__and4b_1
XFILLER_0_119_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07455_ _02018_ _00388_ _03004_ _02040_ VGND VGND VPWR VPWR _04356_ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_826 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10666__A _00819_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07386_ _03576_ _03587_ _03499_ net63 VGND VGND VPWR VPWR _03598_ sky130_fd_sc_hd__and4_1
XFILLER_0_45_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_107 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09125_ _01249_ VGND VGND VPWR VPWR _01250_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_44_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09056_ _01112_ _01174_ VGND VGND VPWR VPWR _01176_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_103_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08007_ _00048_ _00049_ net174 _07048_ VGND VGND VPWR VPWR _00051_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_130_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09958_ _02154_ _02162_ VGND VGND VPWR VPWR _02163_ sky130_fd_sc_hd__nor2_1
X_08909_ _06775_ _00151_ VGND VGND VPWR VPWR _01015_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09889_ _01982_ _01989_ VGND VGND VPWR VPWR _02087_ sky130_fd_sc_hd__or2b_1
X_11920_ _04214_ _04150_ VGND VGND VPWR VPWR _04317_ sky130_fd_sc_hd__and2b_1
XANTENNA__09414__B _00661_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08895__A1 _00508_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07215__A _01284_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11851_ _02663_ _04238_ _04240_ VGND VGND VPWR VPWR _04241_ sky130_fd_sc_hd__and3_1
X_10802_ _03086_ _03087_ VGND VGND VPWR VPWR _03088_ sky130_fd_sc_hd__xnor2_1
X_11782_ _02655_ _02654_ VGND VGND VPWR VPWR _04165_ sky130_fd_sc_hd__or2b_1
XFILLER_0_94_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09430__A _01584_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13521_ _06018_ _03697_ _03699_ _06009_ VGND VGND VPWR VPWR _06060_ sky130_fd_sc_hd__a22o_1
X_10733_ _02885_ _02886_ VGND VGND VPWR VPWR _03012_ sky130_fd_sc_hd__or2_1
XFILLER_0_138_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13452_ _05970_ _05973_ VGND VGND VPWR VPWR _05984_ sky130_fd_sc_hd__or2_1
X_10664_ _02835_ _02837_ VGND VGND VPWR VPWR _02936_ sky130_fd_sc_hd__and2_1
XFILLER_0_82_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12403_ _04839_ _04838_ VGND VGND VPWR VPWR _04848_ sky130_fd_sc_hd__and2b_1
XFILLER_0_3_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09072__A1 _01996_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13383_ _05907_ _05908_ VGND VGND VPWR VPWR _05909_ sky130_fd_sc_hd__or2_1
XFILLER_0_63_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10595_ _00310_ _02855_ _02857_ _00145_ VGND VGND VPWR VPWR _02860_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07885__A _01120_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12334_ _04770_ _04771_ VGND VGND VPWR VPWR _04772_ sky130_fd_sc_hd__and2b_1
XFILLER_0_51_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12265_ _04687_ _04694_ _04695_ VGND VGND VPWR VPWR _04696_ sky130_fd_sc_hd__a21o_1
X_14004_ _06535_ _06545_ _06543_ VGND VGND VPWR VPWR _06591_ sky130_fd_sc_hd__o21ai_1
X_11216_ _03541_ _03542_ VGND VGND VPWR VPWR _03544_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12196_ _03487_ _03512_ _04619_ VGND VGND VPWR VPWR _04621_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_120_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput71 net71 VGND VGND VPWR VPWR prod[15] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_128_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput82 net82 VGND VGND VPWR VPWR prod[25] sky130_fd_sc_hd__clkbuf_4
Xoutput93 net93 VGND VGND VPWR VPWR prod[35] sky130_fd_sc_hd__clkbuf_4
X_11147_ _03458_ _03467_ VGND VGND VPWR VPWR _03468_ sky130_fd_sc_hd__nor2_1
XANTENNA__09127__A2 _01182_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11078_ _03360_ _03355_ _03358_ VGND VGND VPWR VPWR _03392_ sky130_fd_sc_hd__nor3_1
X_10029_ _02152_ _01948_ _01949_ _02240_ VGND VGND VPWR VPWR _02241_ sky130_fd_sc_hd__o31ai_4
XANTENNA__09324__B _00654_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12388__D _01584_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12966__A _05464_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10189__C _00486_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11870__A _06885_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08638__A1 _00439_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13719_ _06270_ _06275_ VGND VGND VPWR VPWR _06278_ sky130_fd_sc_hd__and2b_1
X_07240_ _01000_ VGND VGND VPWR VPWR _01996_ sky130_fd_sc_hd__buf_4
XFILLER_0_144_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__14108__D _02742_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07171_ _00978_ _00705_ _01208_ _00869_ VGND VGND VPWR VPWR _01241_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08810__A1 _00300_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13698__A1 _01289_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08403__B _00460_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13698__B2 _01188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09812_ _02001_ _02002_ VGND VGND VPWR VPWR _02003_ sky130_fd_sc_hd__nor2_2
X_09743_ _01921_ _01926_ VGND VGND VPWR VPWR _01927_ sky130_fd_sc_hd__xor2_1
XANTENNA__07129__A1 net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09674_ _01729_ net143 _01849_ VGND VGND VPWR VPWR _01851_ sky130_fd_sc_hd__nor3_1
XFILLER_0_69_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08625_ _00686_ _00703_ VGND VGND VPWR VPWR _00704_ sky130_fd_sc_hd__xor2_2
XTAP_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12876__A _01504_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08556_ _00599_ _00600_ _00627_ VGND VGND VPWR VPWR _00629_ sky130_fd_sc_hd__and3_1
XTAP_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07507_ _04873_ VGND VGND VPWR VPWR _04928_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_92_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08487_ net182 _00347_ VGND VGND VPWR VPWR _00554_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_848 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10987__A2 _00459_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07438_ _00978_ VGND VGND VPWR VPWR _04169_ sky130_fd_sc_hd__buf_2
XFILLER_0_147_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07369_ _02806_ _03389_ VGND VGND VPWR VPWR _03411_ sky130_fd_sc_hd__or2_4
XFILLER_0_134_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11936__A1 _00004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09108_ _01184_ _01232_ VGND VGND VPWR VPWR _01233_ sky130_fd_sc_hd__xnor2_4
XANTENNA__08016__D net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_767 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10380_ _00486_ _01211_ VGND VGND VPWR VPWR _02625_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_430 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09039_ _01152_ _01154_ _01155_ _01156_ VGND VGND VPWR VPWR _01157_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_103_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_288 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13689__A1 _01289_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12050_ _04137_ _04139_ _04134_ VGND VGND VPWR VPWR _04460_ sky130_fd_sc_hd__a21oi_1
X_11001_ _02971_ _04378_ net47 _00959_ VGND VGND VPWR VPWR _03307_ sky130_fd_sc_hd__and4_1
XANTENNA__12361__B2 _03696_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13592__D _03785_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12952_ _05430_ _05448_ VGND VGND VPWR VPWR _05452_ sky130_fd_sc_hd__and2_1
XFILLER_0_99_255 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11903_ _02335_ _03678_ _04295_ VGND VGND VPWR VPWR _04298_ sky130_fd_sc_hd__a21oi_1
XTAP_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12786__A _01585_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12883_ _05366_ _05375_ VGND VGND VPWR VPWR _05376_ sky130_fd_sc_hd__xor2_1
XTAP_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11834_ _02680_ _04221_ VGND VGND VPWR VPWR _04222_ sky130_fd_sc_hd__xnor2_1
XTAP_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09160__A _01288_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11765_ _02280_ _03682_ VGND VGND VPWR VPWR _04146_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08096__A2 _04895_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10737__C _02758_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_196 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13504_ _06033_ _06039_ VGND VGND VPWR VPWR _06041_ sky130_fd_sc_hd__or2_1
X_10716_ _02890_ _02992_ VGND VGND VPWR VPWR _02994_ sky130_fd_sc_hd__or2_1
X_11696_ _06873_ _01272_ _01211_ _06875_ VGND VGND VPWR VPWR _04071_ sky130_fd_sc_hd__a22o_1
XFILLER_0_83_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10647_ _02895_ _02915_ VGND VGND VPWR VPWR _02918_ sky130_fd_sc_hd__and2_1
X_13435_ _05830_ _05962_ _05965_ VGND VGND VPWR VPWR _05966_ sky130_fd_sc_hd__a21o_1
XFILLER_0_36_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07111__C _00573_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer4 _06142_ VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09596__A2 net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13366_ _05886_ _05889_ VGND VGND VPWR VPWR _05891_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_106_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10578_ _02813_ _02841_ VGND VGND VPWR VPWR _02842_ sky130_fd_sc_hd__xor2_1
XFILLER_0_140_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08504__A net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12317_ _00460_ _02088_ _04749_ VGND VGND VPWR VPWR _04754_ sky130_fd_sc_hd__a21oi_1
X_13297_ _05804_ _05814_ _05819_ VGND VGND VPWR VPWR _05820_ sky130_fd_sc_hd__a21oi_2
X_12248_ _00379_ _03748_ _04677_ VGND VGND VPWR VPWR _04678_ sky130_fd_sc_hd__and3_1
XFILLER_0_139_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12179_ _03589_ _03551_ _03583_ VGND VGND VPWR VPWR _04602_ sky130_fd_sc_hd__a21o_1
XANTENNA__08859__A1 _03587_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08596__D _00258_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08859__B2 _03576_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08410_ _00134_ _00136_ _00287_ _00468_ VGND VGND VPWR VPWR _00469_ sky130_fd_sc_hd__a31o_1
X_09390_ _01539_ _01540_ VGND VGND VPWR VPWR _01541_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08341_ _02138_ _00391_ _00393_ _00344_ VGND VGND VPWR VPWR _00394_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_47_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08272_ _00316_ _00317_ VGND VGND VPWR VPWR _00318_ sky130_fd_sc_hd__nand2_1
XFILLER_0_117_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07223_ _01700_ _01788_ _01799_ VGND VGND VPWR VPWR _01810_ sky130_fd_sc_hd__a21boi_4
XFILLER_0_61_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13368__B1 _02765_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07154_ net1 _01044_ _00923_ net61 VGND VGND VPWR VPWR _01055_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12591__A1 _00745_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12591__B2 _00914_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07085_ net33 VGND VGND VPWR VPWR _00300_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_120_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07675__D _06744_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11692__A1_N _03510_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12343__A1 _01260_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12343__B2 _00755_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07987_ _00028_ _00030_ VGND VGND VPWR VPWR _00031_ sky130_fd_sc_hd__xor2_1
X_09726_ _01681_ _01684_ _01907_ VGND VGND VPWR VPWR _01909_ sky130_fd_sc_hd__a21o_1
XFILLER_0_69_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10657__A1 _00636_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09511__A2 _00459_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09657_ _01829_ _01830_ _01831_ VGND VGND VPWR VPWR _01834_ sky130_fd_sc_hd__a21o_1
XANTENNA__10657__B2 _01156_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08608_ _00668_ _00685_ VGND VGND VPWR VPWR _00686_ sky130_fd_sc_hd__xnor2_2
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09588_ _00991_ _01356_ _01756_ _01757_ _01752_ VGND VGND VPWR VPWR _01758_ sky130_fd_sc_hd__a311o_1
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08539_ _00453_ _02051_ _00458_ _00608_ VGND VGND VPWR VPWR _00610_ sky130_fd_sc_hd__nand4_1
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_848 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11015__A _05181_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11550_ _03907_ _03908_ _03906_ VGND VGND VPWR VPWR _03910_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_147_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10501_ _02754_ _02756_ VGND VGND VPWR VPWR _02757_ sky130_fd_sc_hd__xnor2_1
X_11481_ _03826_ _03832_ _03833_ VGND VGND VPWR VPWR _03834_ sky130_fd_sc_hd__o21a_1
XFILLER_0_107_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13220_ _05744_ _05745_ _05746_ VGND VGND VPWR VPWR _05747_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_107_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10432_ _02680_ _02681_ VGND VGND VPWR VPWR _02682_ sky130_fd_sc_hd__or2_1
XANTENNA__08324__A _00374_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13151_ _05669_ _05670_ VGND VGND VPWR VPWR _05671_ sky130_fd_sc_hd__and2_4
XFILLER_0_20_214 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10363_ _06744_ _03938_ VGND VGND VPWR VPWR _02606_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12102_ _04515_ _04516_ VGND VGND VPWR VPWR _04517_ sky130_fd_sc_hd__nand2_1
XFILLER_0_131_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13082_ _05528_ _05581_ _05582_ _05587_ _05594_ VGND VGND VPWR VPWR _05595_ sky130_fd_sc_hd__o311ai_4
X_10294_ _03268_ _01058_ VGND VGND VPWR VPWR _02530_ sky130_fd_sc_hd__nand2_1
XANTENNA__08538__B1 _00608_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12033_ _04439_ _04440_ VGND VGND VPWR VPWR _04441_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__08994__A _00464_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13984_ _05898_ _05942_ _06567_ VGND VGND VPWR VPWR _06569_ sky130_fd_sc_hd__a21oi_1
X_12935_ _03614_ _05432_ VGND VGND VPWR VPWR _05433_ sky130_fd_sc_hd__xor2_2
XFILLER_0_87_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13405__A _01066_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12866_ _02008_ _02765_ VGND VGND VPWR VPWR _05358_ sky130_fd_sc_hd__nand2_1
XTAP_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07403__A _00322_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11817_ _04185_ _04190_ VGND VGND VPWR VPWR _04204_ sky130_fd_sc_hd__nor2_1
XTAP_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12797_ _00914_ _01933_ _05101_ _05281_ VGND VGND VPWR VPWR _05282_ sky130_fd_sc_hd__a31o_1
XTAP_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12270__B1 _01250_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07816__A2 net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11748_ _02616_ _02633_ VGND VGND VPWR VPWR _04128_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09018__A1 _03543_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11679_ _04049_ _04050_ _04042_ _04044_ VGND VGND VPWR VPWR _04052_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_71_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13418_ _05946_ _05947_ VGND VGND VPWR VPWR _05948_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13349_ _01600_ _01585_ _02306_ _02857_ VGND VGND VPWR VPWR _05872_ sky130_fd_sc_hd__nand4_1
XFILLER_0_11_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10584__B1 _02305_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12325__A1 _01289_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07910_ _06932_ _06934_ _07038_ VGND VGND VPWR VPWR _07039_ sky130_fd_sc_hd__a21o_1
X_08890_ _06966_ _04906_ _04928_ _06965_ VGND VGND VPWR VPWR _00994_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07841_ _06963_ _06967_ _06968_ _06969_ VGND VGND VPWR VPWR _06970_ sky130_fd_sc_hd__or4_1
XANTENNA__12203__B _04627_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07772_ _01208_ _04851_ net4 _00705_ VGND VGND VPWR VPWR _06901_ sky130_fd_sc_hd__a22o_1
XANTENNA__13018__C _05524_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09511_ _06494_ _00459_ _01671_ VGND VGND VPWR VPWR _01673_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_78_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09442_ _06439_ _00414_ _00574_ _02018_ VGND VGND VPWR VPWR _01598_ sky130_fd_sc_hd__a22o_1
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09373_ _01388_ _01391_ _01521_ VGND VGND VPWR VPWR _01522_ sky130_fd_sc_hd__o21a_1
XFILLER_0_59_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08324_ _00374_ VGND VGND VPWR VPWR _00375_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__13969__B _06552_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12873__B _03748_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08255_ _00157_ _00159_ _00144_ _00298_ VGND VGND VPWR VPWR _00299_ sky130_fd_sc_hd__and4_1
XANTENNA__07967__B _01120_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10674__A _00294_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_531 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07206_ _01580_ _01613_ VGND VGND VPWR VPWR _01624_ sky130_fd_sc_hd__or2b_1
XFILLER_0_131_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08186_ _00228_ _00226_ VGND VGND VPWR VPWR _00230_ sky130_fd_sc_hd__and2b_1
XFILLER_0_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10824__D net57 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07137_ net23 VGND VGND VPWR VPWR _00869_ sky130_fd_sc_hd__buf_8
XFILLER_0_113_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11001__C net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09709_ _01682_ _01683_ VGND VGND VPWR VPWR _01890_ sky130_fd_sc_hd__nor2_1
X_10981_ _03283_ _03284_ VGND VGND VPWR VPWR _03285_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09496__A1 _01284_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10849__A _05742_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12720_ _04993_ _05031_ VGND VGND VPWR VPWR _05197_ sky130_fd_sc_hd__xor2_1
XFILLER_0_97_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09422__B _00745_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08319__A _00354_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12651_ _05120_ _05080_ VGND VGND VPWR VPWR _05121_ sky130_fd_sc_hd__xnor2_1
X_11602_ _03961_ _03963_ VGND VGND VPWR VPWR _03967_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12582_ _05043_ _05044_ VGND VGND VPWR VPWR _05045_ sky130_fd_sc_hd__or2b_1
XFILLER_0_25_306 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11533_ _03886_ _03890_ VGND VGND VPWR VPWR _03891_ sky130_fd_sc_hd__xor2_2
XANTENNA__13598__C _01250_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_434 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09795__D _01586_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11464_ _00497_ _03681_ VGND VGND VPWR VPWR _03815_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13203_ _05455_ _05726_ _05727_ VGND VGND VPWR VPWR _05728_ sky130_fd_sc_hd__o21ai_2
X_10415_ _02646_ _02442_ _02647_ _02662_ VGND VGND VPWR VPWR _02663_ sky130_fd_sc_hd__or4_2
X_14183_ _06750_ _06782_ _06769_ VGND VGND VPWR VPWR _06783_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_104_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11395_ _03736_ _03737_ _06765_ _03738_ VGND VGND VPWR VPWR _03739_ sky130_fd_sc_hd__and4bb_1
X_10346_ _02583_ _02586_ VGND VGND VPWR VPWR _02588_ sky130_fd_sc_hd__xnor2_2
X_13134_ _05649_ _05651_ VGND VGND VPWR VPWR _05652_ sky130_fd_sc_hd__nor2_2
XFILLER_0_131_591 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13065_ _05565_ _05567_ VGND VGND VPWR VPWR _05576_ sky130_fd_sc_hd__xor2_2
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10277_ _02509_ _02511_ VGND VGND VPWR VPWR _02512_ sky130_fd_sc_hd__xor2_1
XFILLER_0_29_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12016_ _04421_ _04346_ VGND VGND VPWR VPWR _04423_ sky130_fd_sc_hd__or2_1
XFILLER_0_136_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08220__C _00262_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap2 net180 VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13967_ _06471_ _06473_ _06474_ VGND VGND VPWR VPWR _06551_ sky130_fd_sc_hd__nand3_1
X_12918_ _01108_ _01183_ VGND VGND VPWR VPWR _05415_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13898_ _06471_ _06473_ _06474_ VGND VGND VPWR VPWR _06475_ sky130_fd_sc_hd__a21o_1
XFILLER_0_88_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12849_ _01585_ _01060_ _05268_ VGND VGND VPWR VPWR _05339_ sky130_fd_sc_hd__and3_1
XFILLER_0_29_634 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10178__A1_N _06744_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08040_ _00081_ _00082_ _07077_ VGND VGND VPWR VPWR _00084_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_126_385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12546__A1 _00393_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_142_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12546__B2 _00390_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09991_ _01535_ _01676_ _01902_ _01900_ VGND VGND VPWR VPWR _02199_ sky130_fd_sc_hd__a31o_1
XFILLER_0_12_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08942_ _00765_ _00887_ _00886_ VGND VGND VPWR VPWR _01051_ sky130_fd_sc_hd__a21o_1
XANTENNA__09507__B _00607_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09714__A2 _00608_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08873_ _00971_ _00974_ VGND VGND VPWR VPWR _00975_ sky130_fd_sc_hd__xor2_1
XFILLER_0_36_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07824_ _00420_ net39 net38 net177 VGND VGND VPWR VPWR _06953_ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07755_ _02259_ _00508_ VGND VGND VPWR VPWR _06884_ sky130_fd_sc_hd__nand2_2
X_07686_ net26 net64 VGND VGND VPWR VPWR _06815_ sky130_fd_sc_hd__nand2_1
XANTENNA__12482__B1 _03762_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09425_ _01574_ _01267_ _01578_ VGND VGND VPWR VPWR _01579_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_137_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09356_ _01369_ VGND VGND VPWR VPWR _01504_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__12234__B1 _01248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12785__A1 _01586_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08307_ _00089_ _00090_ VGND VGND VPWR VPWR _00357_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09287_ _01112_ _01174_ VGND VGND VPWR VPWR _01429_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08238_ _00280_ _00281_ VGND VGND VPWR VPWR _00282_ sky130_fd_sc_hd__or2_1
XFILLER_0_90_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08169_ _06120_ _00212_ _06153_ VGND VGND VPWR VPWR _00213_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10548__B1 _02730_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10200_ _06450_ _02427_ VGND VGND VPWR VPWR _02428_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11180_ _03500_ _03501_ _03502_ _03503_ VGND VGND VPWR VPWR _03504_ sky130_fd_sc_hd__nor4_1
XFILLER_0_113_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10851__B _03268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10131_ _00151_ _01517_ _02351_ VGND VGND VPWR VPWR _02352_ sky130_fd_sc_hd__and3_1
X_10062_ _01646_ _01643_ _01837_ _02045_ _02276_ VGND VGND VPWR VPWR _02277_ sky130_fd_sc_hd__a41o_1
XANTENNA__07218__A _00442_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13821_ _04714_ _03683_ VGND VGND VPWR VPWR _06390_ sky130_fd_sc_hd__nand2_1
XANTENNA__09433__A _00157_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10579__A _00143_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13265__A2 _05524_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13752_ _06312_ _06313_ VGND VGND VPWR VPWR _06314_ sky130_fd_sc_hd__nor2_1
X_10964_ _03261_ _03264_ VGND VGND VPWR VPWR _03266_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12703_ _04690_ _04691_ VGND VGND VPWR VPWR _05178_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_97_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13683_ _06116_ _06237_ VGND VGND VPWR VPWR _06238_ sky130_fd_sc_hd__xnor2_4
XANTENNA__12794__A _00914_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10895_ _03185_ _03184_ VGND VGND VPWR VPWR _03190_ sky130_fd_sc_hd__and2b_1
X_12634_ _02168_ _05100_ _05101_ VGND VGND VPWR VPWR _05102_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_31_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_423 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12565_ _05012_ _05025_ VGND VGND VPWR VPWR _05026_ sky130_fd_sc_hd__xor2_2
XFILLER_0_80_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11516_ _03853_ _03856_ VGND VGND VPWR VPWR _03873_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__07400__B _00322_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12496_ _04948_ _04949_ VGND VGND VPWR VPWR _04951_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_124_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08215__C _00257_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11447_ _03793_ _03794_ _03796_ VGND VGND VPWR VPWR _03797_ sky130_fd_sc_hd__and3_1
XANTENNA__10003__A2 _04037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09608__A _01585_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14166_ _06764_ _06741_ VGND VGND VPWR VPWR _06766_ sky130_fd_sc_hd__or2_1
X_11378_ _03717_ _03720_ VGND VGND VPWR VPWR _03721_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10329_ _02567_ _02568_ VGND VGND VPWR VPWR _02569_ sky130_fd_sc_hd__xor2_1
X_13117_ _03669_ _05633_ VGND VGND VPWR VPWR _05634_ sky130_fd_sc_hd__xnor2_2
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14097_ _06684_ _06692_ VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__xor2_4
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08231__B _06775_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13048_ _00376_ _00391_ _00393_ _00381_ VGND VGND VPWR VPWR _05558_ sky130_fd_sc_hd__a22oi_2
XANTENNA__12969__A _05455_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08904__B1 _00114_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10489__A _01473_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07540_ _05082_ _05280_ VGND VGND VPWR VPWR _05291_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_89_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07471_ _04488_ _04499_ _04521_ VGND VGND VPWR VPWR _04532_ sky130_fd_sc_hd__and3_2
XFILLER_0_76_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09880__A1 _03554_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09880__B2 _00508_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09210_ _01329_ _01343_ VGND VGND VPWR VPWR _01344_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12216__B1 _01249_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_626 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09141_ _01257_ _01202_ _01266_ VGND VGND VPWR VPWR _01268_ sky130_fd_sc_hd__and3_1
XFILLER_0_146_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_650 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13312__B _05833_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09072_ _01996_ _03894_ _00920_ _00919_ VGND VGND VPWR VPWR _01193_ sky130_fd_sc_hd__a31o_1
XFILLER_0_115_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08023_ _06909_ _07066_ _07065_ VGND VGND VPWR VPWR _00067_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_114_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11767__B _02335_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09974_ _02153_ _02179_ VGND VGND VPWR VPWR _02180_ sky130_fd_sc_hd__or2_2
XANTENNA__07683__D net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08925_ _01030_ _01031_ VGND VGND VPWR VPWR _01032_ sky130_fd_sc_hd__or2_2
X_08856_ _00954_ _00955_ VGND VGND VPWR VPWR _00957_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__12598__B _03740_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07807_ _06658_ _06669_ VGND VGND VPWR VPWR _06936_ sky130_fd_sc_hd__and2_1
X_08787_ _00707_ _00709_ VGND VGND VPWR VPWR _00882_ sky130_fd_sc_hd__nor2_1
X_07738_ _06865_ _06866_ VGND VGND VPWR VPWR _06867_ sky130_fd_sc_hd__and2b_1
XANTENNA__11007__B _01664_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07669_ _06142_ _06175_ _06406_ _06615_ _06680_ VGND VGND VPWR VPWR _06691_ sky130_fd_sc_hd__a2111oi_4
XANTENNA__07204__C _01208_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09408_ _01559_ _01487_ _01490_ VGND VGND VPWR VPWR _01561_ sky130_fd_sc_hd__and3_1
XANTENNA__07882__B1 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10680_ _00366_ _02982_ _01546_ _02156_ VGND VGND VPWR VPWR _02954_ sky130_fd_sc_hd__and4_1
XFILLER_0_47_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12758__A1 _00457_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07501__A _04851_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09339_ _01445_ _01446_ _01483_ VGND VGND VPWR VPWR _01485_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_35_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12350_ _04788_ _04789_ VGND VGND VPWR VPWR _04790_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11301_ _03634_ _03636_ VGND VGND VPWR VPWR _03637_ sky130_fd_sc_hd__and2_1
XANTENNA__11958__A _00138_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12281_ _01066_ VGND VGND VPWR VPWR _04714_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_105_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14020_ _06492_ _06507_ _06607_ _06608_ _06240_ VGND VGND VPWR VPWR _06609_ sky130_fd_sc_hd__o32a_2
X_11232_ _03556_ _03559_ VGND VGND VPWR VPWR _03561_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08332__A _00383_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11163_ _03461_ _03462_ VGND VGND VPWR VPWR _03485_ sky130_fd_sc_hd__xnor2_2
XANTENNA__09147__B _01405_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11396__C _01254_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10114_ _02301_ _02332_ VGND VGND VPWR VPWR _02333_ sky130_fd_sc_hd__xnor2_2
X_11094_ _03406_ _03408_ VGND VGND VPWR VPWR _03409_ sky130_fd_sc_hd__nand2_1
XANTENNA__07890__B _00475_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10045_ _02256_ _02257_ VGND VGND VPWR VPWR _02258_ sky130_fd_sc_hd__nor2_1
XANTENNA__12004__D _01780_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_output126_A net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13804_ _02190_ _03684_ _03680_ _02188_ VGND VGND VPWR VPWR _06371_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_98_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11996_ _04328_ _04398_ _04399_ VGND VGND VPWR VPWR _04401_ sky130_fd_sc_hd__and3_1
XFILLER_0_86_824 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13735_ _00916_ _02730_ _06294_ VGND VGND VPWR VPWR _06295_ sky130_fd_sc_hd__and3_1
X_10947_ _03189_ _03205_ _03242_ _03245_ _03247_ VGND VGND VPWR VPWR _03248_ sky130_fd_sc_hd__a41o_1
XANTENNA__09862__A1 _00519_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__09610__B _01780_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13666_ _06217_ _06218_ VGND VGND VPWR VPWR _06220_ sky130_fd_sc_hd__nand2_2
XFILLER_0_38_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10878_ _03168_ _03171_ VGND VGND VPWR VPWR _03172_ sky130_fd_sc_hd__and2_1
XANTENNA__08507__A _00574_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12617_ _05059_ _05083_ VGND VGND VPWR VPWR _05084_ sky130_fd_sc_hd__xor2_1
X_13597_ _01413_ _01249_ _02856_ _01180_ VGND VGND VPWR VPWR _06144_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07130__B net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12548_ _05007_ _04954_ VGND VGND VPWR VPWR _05008_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12479_ _04919_ _04931_ VGND VGND VPWR VPWR _04932_ sky130_fd_sc_hd__and2_1
XFILLER_0_112_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14218_ _00464_ _00344_ VGND VGND VPWR VPWR _06804_ sky130_fd_sc_hd__and2_1
XANTENNA__09917__A2 _02117_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14149_ _06746_ _06729_ VGND VGND VPWR VPWR _06748_ sky130_fd_sc_hd__or2b_1
XTAP_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13477__A2 _01956_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08710_ _00790_ _00796_ VGND VGND VPWR VPWR _00797_ sky130_fd_sc_hd__and2_1
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09690_ _04939_ _00379_ VGND VGND VPWR VPWR _01869_ sky130_fd_sc_hd__nand2_1
XANTENNA__12685__B1 _05150_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09073__A _05445_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08641_ _00718_ _00719_ VGND VGND VPWR VPWR _00722_ sky130_fd_sc_hd__xor2_1
Xrebuffer14 _00588_ VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__buf_1
XANTENNA__12211__B _00379_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xrebuffer25 _07061_ VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__clkbuf_1
Xrebuffer36 _05967_ VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_89_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08572_ _00644_ _00645_ VGND VGND VPWR VPWR _00646_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07523_ _03147_ _00355_ _02960_ net60 VGND VGND VPWR VPWR _05104_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07454_ _01996_ _00901_ _00366_ _02982_ VGND VGND VPWR VPWR _04345_ sky130_fd_sc_hd__nand4_2
XFILLER_0_92_838 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10666__B _00818_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07385_ _00978_ VGND VGND VPWR VPWR _03587_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_146_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09124_ _01248_ VGND VGND VPWR VPWR _01249_ sky130_fd_sc_hd__buf_4
XFILLER_0_115_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09055_ _01166_ _01173_ VGND VGND VPWR VPWR _01174_ sky130_fd_sc_hd__xor2_2
XFILLER_0_115_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_651 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08006_ _07047_ _07048_ _00048_ _00049_ VGND VGND VPWR VPWR _00050_ sky130_fd_sc_hd__o211a_1
XFILLER_0_130_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09957_ _02155_ _02161_ VGND VGND VPWR VPWR _02162_ sky130_fd_sc_hd__xnor2_1
X_08908_ _06775_ _00095_ _00826_ _00656_ _00258_ VGND VGND VPWR VPWR _01014_ sky130_fd_sc_hd__a32o_1
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09888_ _02085_ VGND VGND VPWR VPWR _02086_ sky130_fd_sc_hd__inv_2
X_08839_ _00751_ _00761_ VGND VGND VPWR VPWR _00938_ sky130_fd_sc_hd__nand2_1
XANTENNA__09414__C net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08895__A2 _00158_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11850_ _04223_ _04239_ VGND VGND VPWR VPWR _04240_ sky130_fd_sc_hd__nor2_1
XANTENNA__07215__B _00300_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10801_ _06483_ _01933_ VGND VGND VPWR VPWR _03087_ sky130_fd_sc_hd__nand2_1
XFILLER_0_138_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11781_ _04157_ _04163_ VGND VGND VPWR VPWR _04164_ sky130_fd_sc_hd__xor2_1
XFILLER_0_95_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13520_ _06057_ _06058_ VGND VGND VPWR VPWR _06059_ sky130_fd_sc_hd__nor2_1
X_10732_ _03008_ _03010_ VGND VGND VPWR VPWR _03011_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08327__A _00378_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13451_ _05981_ _05982_ VGND VGND VPWR VPWR _05983_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10663_ _02930_ _02934_ VGND VGND VPWR VPWR _02935_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_82_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12402_ _04841_ _04844_ _04846_ VGND VGND VPWR VPWR _04847_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_35_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10594_ _00145_ _00310_ _02856_ _02858_ VGND VGND VPWR VPWR _02859_ sky130_fd_sc_hd__nand4_1
X_13382_ _05900_ _05906_ VGND VGND VPWR VPWR _05908_ sky130_fd_sc_hd__nor2_1
XANTENNA__09072__A2 _03894_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_130 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12333_ _04744_ _04746_ VGND VGND VPWR VPWR _04771_ sky130_fd_sc_hd__xor2_1
XANTENNA__07885__B net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10592__A _02305_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12264_ _04678_ _04684_ _04685_ VGND VGND VPWR VPWR _04695_ sky130_fd_sc_hd__o21a_1
XFILLER_0_50_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14003_ _06588_ _06589_ VGND VGND VPWR VPWR _06590_ sky130_fd_sc_hd__and2_1
X_11215_ _03539_ _03540_ VGND VGND VPWR VPWR _03542_ sky130_fd_sc_hd__nor2_1
X_12195_ _03484_ _03486_ VGND VGND VPWR VPWR _04619_ sky130_fd_sc_hd__or2_1
Xoutput72 net72 VGND VGND VPWR VPWR prod[16] sky130_fd_sc_hd__clkbuf_4
Xoutput83 net83 VGND VGND VPWR VPWR prod[26] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11146_ _03461_ _03462_ _03465_ VGND VGND VPWR VPWR _03467_ sky130_fd_sc_hd__o21ai_2
Xoutput94 net94 VGND VGND VPWR VPWR prod[36] sky130_fd_sc_hd__buf_2
X_11077_ _03331_ _03390_ VGND VGND VPWR VPWR _03391_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12312__A _00415_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10028_ _02236_ _02239_ VGND VGND VPWR VPWR _02240_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_144_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_312 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11870__B _01780_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11979_ _04380_ _04381_ VGND VGND VPWR VPWR _04382_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13718_ _06268_ _06276_ VGND VGND VPWR VPWR _06277_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_827 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07141__A _00891_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13649_ _06191_ _06195_ _06200_ VGND VGND VPWR VPWR _06201_ sky130_fd_sc_hd__and3_1
XFILLER_0_144_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07170_ net26 VGND VGND VPWR VPWR _01230_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__08810__A2 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09068__A _02456_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13698__A2 _02726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09811_ _01998_ _02000_ VGND VGND VPWR VPWR _02002_ sky130_fd_sc_hd__and2_1
XANTENNA__08700__A _01350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09742_ _01924_ _01925_ VGND VGND VPWR VPWR _01926_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07129__A2 net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09673_ _01729_ net143 _01849_ VGND VGND VPWR VPWR _01850_ sky130_fd_sc_hd__o21a_1
XFILLER_0_118_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08624_ _00687_ _00702_ VGND VGND VPWR VPWR _00703_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_77_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12876__B _01249_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08555_ _00603_ _00626_ VGND VGND VPWR VPWR _00627_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10677__A _05181_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13053__A _05546_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07506_ _04906_ VGND VGND VPWR VPWR _04917_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_119_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08486_ _00550_ _00551_ VGND VGND VPWR VPWR _00553_ sky130_fd_sc_hd__or2_1
XFILLER_0_64_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12830__B1 _04600_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07437_ _04070_ _04147_ VGND VGND VPWR VPWR _04158_ sky130_fd_sc_hd__nand2_1
XANTENNA__09039__C1 _01156_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12892__A _00784_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07368_ _02806_ _03389_ VGND VGND VPWR VPWR _03400_ sky130_fd_sc_hd__and2_4
XANTENNA__11397__B1 _02119_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09107_ _01229_ _01231_ VGND VGND VPWR VPWR _01232_ sky130_fd_sc_hd__or2b_2
XANTENNA__11936__A2 _01585_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07299_ _00792_ _00781_ VGND VGND VPWR VPWR _02642_ sky130_fd_sc_hd__or2b_1
XFILLER_0_32_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09038_ _00526_ VGND VGND VPWR VPWR _01156_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_60_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13689__A2 _02730_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_486 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11000_ _04378_ net47 _00959_ _02971_ VGND VGND VPWR VPWR _03306_ sky130_fd_sc_hd__a22o_1
XANTENNA__12361__A2 _00604_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12951_ _05018_ _05450_ VGND VGND VPWR VPWR _05451_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_99_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11902_ _03070_ _03682_ _04292_ _04293_ VGND VGND VPWR VPWR _04297_ sky130_fd_sc_hd__o2bb2a_1
XTAP_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__11872__A1 _07004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12882_ _05367_ _05374_ VGND VGND VPWR VPWR _05375_ sky130_fd_sc_hd__xor2_1
XTAP_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12786__B _01059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09441__A _06439_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11833_ _04220_ _04188_ VGND VGND VPWR VPWR _04221_ sky130_fd_sc_hd__nor2_1
XTAP_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11764_ _02135_ _04143_ _04144_ VGND VGND VPWR VPWR _04145_ sky130_fd_sc_hd__a21bo_1
XANTENNA__08057__A net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13503_ _06033_ _06039_ VGND VGND VPWR VPWR _06040_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10737__D _02721_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10715_ _02887_ _02889_ VGND VGND VPWR VPWR _02992_ sky130_fd_sc_hd__and2_1
XFILLER_0_83_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11695_ _06964_ _06875_ _01272_ _01211_ VGND VGND VPWR VPWR _04069_ sky130_fd_sc_hd__nand4_1
XFILLER_0_71_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13377__A1 _01504_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07896__A _02719_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13377__B2 _01508_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13434_ _05846_ _05961_ _05964_ VGND VGND VPWR VPWR _05965_ sky130_fd_sc_hd__a21o_1
X_10646_ _02895_ _02915_ VGND VGND VPWR VPWR _02917_ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07111__D net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer5 _05522_ VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__buf_1
XFILLER_0_3_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13365_ _02765_ _05887_ _05888_ VGND VGND VPWR VPWR _05889_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_134_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10577_ _02830_ _02838_ _02840_ VGND VGND VPWR VPWR _02841_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_779 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__13824__A2_N _03683_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12316_ _04739_ _04751_ VGND VGND VPWR VPWR _04753_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13296_ _05739_ _05734_ _05817_ VGND VGND VPWR VPWR _05819_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_121_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12247_ _00378_ _02119_ _04674_ _04676_ VGND VGND VPWR VPWR _04677_ sky130_fd_sc_hd__a31o_1
XANTENNA_output70_A net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12178_ _03677_ _04600_ VGND VGND VPWR VPWR _04601_ sky130_fd_sc_hd__xor2_2
XFILLER_0_48_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11129_ _03261_ _03264_ _03300_ _03303_ _03262_ VGND VGND VPWR VPWR _03448_ sky130_fd_sc_hd__a311o_1
XFILLER_0_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08859__A2 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08340_ _00392_ VGND VGND VPWR VPWR _00393_ sky130_fd_sc_hd__buf_4
XFILLER_0_46_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08271_ _00148_ _00315_ VGND VGND VPWR VPWR _00317_ sky130_fd_sc_hd__or2_1
XFILLER_0_144_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07222_ _01624_ _01678_ _01689_ VGND VGND VPWR VPWR _01799_ sky130_fd_sc_hd__a21o_1
XANTENNA__13368__B2 _02008_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07153_ net62 VGND VGND VPWR VPWR _01044_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_144_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__14135__C _02742_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12591__A2 _02855_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10960__A _00145_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07986_ _06949_ _07028_ _00029_ VGND VGND VPWR VPWR _00030_ sky130_fd_sc_hd__a21oi_1
X_09725_ _01681_ _01684_ _01680_ VGND VGND VPWR VPWR _01907_ sky130_fd_sc_hd__o21a_1
XFILLER_0_97_705 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09656_ _01829_ _01830_ _01831_ VGND VGND VPWR VPWR _01833_ sky130_fd_sc_hd__nand3_4
XANTENNA__10657__A2 _02765_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09261__A _00608_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08607_ _00484_ _00684_ VGND VGND VPWR VPWR _00685_ sky130_fd_sc_hd__xnor2_2
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09587_ _01354_ _01486_ _01756_ _01357_ VGND VGND VPWR VPWR _01757_ sky130_fd_sc_hd__a2bb2o_1
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08538_ _02051_ _00458_ _00608_ _00442_ VGND VGND VPWR VPWR _00609_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10200__A _06450_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_186 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11015__B net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08469_ _00532_ _00533_ VGND VGND VPWR VPWR _00534_ sky130_fd_sc_hd__and2b_1
XFILLER_0_37_359 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10500_ _02741_ _02755_ VGND VGND VPWR VPWR _02756_ sky130_fd_sc_hd__nor2_1
XFILLER_0_135_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11480_ _03823_ _03825_ VGND VGND VPWR VPWR _03833_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10431_ _02466_ _02679_ VGND VGND VPWR VPWR _02681_ sky130_fd_sc_hd__and2_1
X_13150_ _04025_ _04595_ VGND VGND VPWR VPWR _05670_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_21_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10362_ _06744_ _03894_ _02400_ _02403_ VGND VGND VPWR VPWR _02605_ sky130_fd_sc_hd__a31o_1
XFILLER_0_115_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12101_ _04427_ _04447_ VGND VGND VPWR VPWR _04516_ sky130_fd_sc_hd__nand2_1
XANTENNA__11790__B1 net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13081_ _05563_ _05589_ _05591_ _05593_ VGND VGND VPWR VPWR _05594_ sky130_fd_sc_hd__a31oi_2
X_10293_ _05577_ net49 _02326_ _02323_ VGND VGND VPWR VPWR _02529_ sky130_fd_sc_hd__a31o_1
XFILLER_0_130_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__08538__A1 _02051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12032_ _04438_ _04428_ VGND VGND VPWR VPWR _04440_ sky130_fd_sc_hd__and2b_1
XANTENNA__08538__B2 _00442_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08340__A _00392_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13983_ _05898_ _05942_ _06567_ VGND VGND VPWR VPWR _06568_ sky130_fd_sc_hd__and3_1
XANTENNA__08994__B _01062_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12934_ _05431_ _03612_ _03619_ VGND VGND VPWR VPWR _05432_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_34_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07933__A2_N net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13405__B _03414_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12865_ _05353_ _05355_ VGND VGND VPWR VPWR _05356_ sky130_fd_sc_hd__xor2_1
XTAP_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_805 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07403__B _03773_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11816_ _04172_ _04177_ _04184_ VGND VGND VPWR VPWR _04203_ sky130_fd_sc_hd__and3_1
XTAP_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12796_ _00389_ _00392_ _02168_ _02723_ VGND VGND VPWR VPWR _05281_ sky130_fd_sc_hd__and4_1
XTAP_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11747_ _04126_ VGND VGND VPWR VPWR _04127_ sky130_fd_sc_hd__inv_2
XANTENNA__12270__A1 _03414_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12270__B2 _01066_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09018__A2 _00144_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11678_ _04042_ _04044_ _04049_ _04050_ VGND VGND VPWR VPWR _04051_ sky130_fd_sc_hd__o211a_1
XFILLER_0_126_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13417_ _05943_ _05944_ _05853_ VGND VGND VPWR VPWR _05947_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08226__B1 _00268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10629_ _00819_ _02735_ VGND VGND VPWR VPWR _02898_ sky130_fd_sc_hd__nand2_1
XFILLER_0_113_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13348_ _01584_ _02306_ _02305_ _01586_ VGND VGND VPWR VPWR _05871_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10584__A1 _04895_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10584__B2 _04928_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13279_ _05793_ _05801_ VGND VGND VPWR VPWR _05802_ sky130_fd_sc_hd__and2_1
XFILLER_0_121_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_782 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08250__A _00151_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07840_ _06878_ _06879_ VGND VGND VPWR VPWR _06969_ sky130_fd_sc_hd__and2b_1
XFILLER_0_75_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07771_ _00705_ _00573_ _04851_ net4 VGND VGND VPWR VPWR _06900_ sky130_fd_sc_hd__and4_1
X_09510_ _06494_ _00458_ _01671_ VGND VGND VPWR VPWR _01672_ sky130_fd_sc_hd__and3_1
XFILLER_0_79_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09441_ _06439_ _02018_ _00574_ VGND VGND VPWR VPWR _01597_ sky130_fd_sc_hd__and3_1
XFILLER_0_93_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09372_ _01516_ _01520_ VGND VGND VPWR VPWR _01521_ sky130_fd_sc_hd__xor2_1
XFILLER_0_47_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09584__B_N _01752_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08323_ _00373_ VGND VGND VPWR VPWR _00374_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_145_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08254_ _00158_ VGND VGND VPWR VPWR _00298_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_145_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07967__C _07010_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10674__B _02857_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07205_ _01076_ net33 _01591_ _01602_ VGND VGND VPWR VPWR _01613_ sky130_fd_sc_hd__a31o_1
XFILLER_0_15_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08185_ _00226_ _00228_ VGND VGND VPWR VPWR _00229_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_131_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__09965__B1 _02169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07136_ _00847_ VGND VGND VPWR VPWR _00858_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11001__D _00959_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10327__A1 _00613_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__14069__A2 _02743_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07969_ _00009_ _00012_ VGND VGND VPWR VPWR _00013_ sky130_fd_sc_hd__xor2_1
X_09708_ _01869_ _01888_ VGND VGND VPWR VPWR _01889_ sky130_fd_sc_hd__xor2_2
X_10980_ _00158_ _00457_ VGND VGND VPWR VPWR _03284_ sky130_fd_sc_hd__nand2_1
XANTENNA__09496__A2 net49 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10849__B _00541_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07504__A _04862_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09639_ _00300_ net19 _01565_ _01567_ VGND VGND VPWR VPWR _01814_ sky130_fd_sc_hd__a31o_1
XFILLER_0_38_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12650_ _05081_ _05073_ VGND VGND VPWR VPWR _05120_ sky130_fd_sc_hd__or2b_1
XFILLER_0_77_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11601_ _03830_ _03965_ VGND VGND VPWR VPWR _03966_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12581_ _00742_ _02849_ _02304_ _00392_ VGND VGND VPWR VPWR _05044_ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11532_ _03887_ _03884_ VGND VGND VPWR VPWR _03890_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_556 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11463_ _03812_ _03813_ VGND VGND VPWR VPWR _03814_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13202_ _05457_ _05469_ VGND VGND VPWR VPWR _05727_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10414_ _02660_ _02661_ VGND VGND VPWR VPWR _02662_ sky130_fd_sc_hd__nor2_1
X_14182_ _06770_ VGND VGND VPWR VPWR _06782_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11394_ _02119_ VGND VGND VPWR VPWR _03738_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_60_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11763__B1 _02134_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13133_ _05635_ _05650_ VGND VGND VPWR VPWR _05651_ sky130_fd_sc_hd__or2b_4
X_10345_ _02584_ _02377_ _02585_ VGND VGND VPWR VPWR _02586_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_103_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13064_ _05573_ _05574_ VGND VGND VPWR VPWR _05575_ sky130_fd_sc_hd__nor2_2
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10276_ _04081_ net54 VGND VGND VPWR VPWR _02511_ sky130_fd_sc_hd__nand2_1
XANTENNA__08070__A _00101_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12015_ _04419_ _04420_ VGND VGND VPWR VPWR _04421_ sky130_fd_sc_hd__nor2_1
XANTENNA__10105__A _00628_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07195__B1 _01208_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08220__D _00263_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13966_ _06352_ _06548_ VGND VGND VPWR VPWR _06550_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07414__A _02127_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13135__B _05636_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12917_ _05411_ _05413_ VGND VGND VPWR VPWR _05414_ sky130_fd_sc_hd__or2b_1
XFILLER_0_76_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12491__A1 _00613_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13897_ _06468_ _06469_ VGND VGND VPWR VPWR _06474_ sky130_fd_sc_hd__xor2_1
XANTENNA__12491__B2 _00612_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10145__A2_N _04048_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12848_ _05268_ _05270_ VGND VGND VPWR VPWR _05338_ sky130_fd_sc_hd__or2b_1
XTAP_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12779_ _04728_ _04732_ _04735_ _04729_ VGND VGND VPWR VPWR _05262_ sky130_fd_sc_hd__a31o_1
XTAP_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12546__A2 _00459_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09947__B1 _02150_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09990_ _02185_ _02197_ VGND VGND VPWR VPWR _02198_ sky130_fd_sc_hd__xnor2_1
X_08941_ _00943_ _01049_ VGND VGND VPWR VPWR _01050_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_110_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08872_ _00615_ _00972_ _00973_ VGND VGND VPWR VPWR _00974_ sky130_fd_sc_hd__and3_1
XANTENNA__10015__A _00459_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07823_ _00420_ net177 net39 net38 VGND VGND VPWR VPWR _06952_ sky130_fd_sc_hd__and4_1
XFILLER_0_29_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07754_ _06856_ _06882_ VGND VGND VPWR VPWR _06883_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11772__C _01996_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12230__A _01517_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07685_ _06812_ _06813_ VGND VGND VPWR VPWR _06814_ sky130_fd_sc_hd__and2b_1
XFILLER_0_67_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12482__B2 _00612_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09424_ _01576_ _01577_ VGND VGND VPWR VPWR _01578_ sky130_fd_sc_hd__and2_1
XFILLER_0_94_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09355_ _01367_ _01373_ VGND VGND VPWR VPWR _01502_ sky130_fd_sc_hd__nor2_1
XANTENNA__12234__A1 _00778_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12234__B2 _00783_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13699__C _02427_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_136_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13061__A _05559_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08306_ _06985_ _07082_ VGND VGND VPWR VPWR _00356_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12785__A2 _01059_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09286_ _01309_ _01426_ VGND VGND VPWR VPWR _01428_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_145_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08237_ _00108_ _00279_ VGND VGND VPWR VPWR _00281_ sky130_fd_sc_hd__and2_1
XFILLER_0_62_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08168_ _02445_ _02883_ _03477_ net140 VGND VGND VPWR VPWR _00212_ sky130_fd_sc_hd__a31o_1
XFILLER_0_43_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10548__A1 _00818_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10548__B2 _00819_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07119_ _00661_ VGND VGND VPWR VPWR _00672_ sky130_fd_sc_hd__buf_4
X_08099_ _00142_ VGND VGND VPWR VPWR _00143_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_30_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10130_ _00094_ _00784_ VGND VGND VPWR VPWR _02351_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10061_ _01833_ _01835_ _02044_ VGND VGND VPWR VPWR _02276_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07218__B _00989_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13820_ _01955_ _06387_ _06388_ VGND VGND VPWR VPWR _06389_ sky130_fd_sc_hd__a21bo_1
XANTENNA__09433__B _01585_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13265__A3 _05593_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10579__B _04906_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13751_ _06309_ _06310_ VGND VGND VPWR VPWR _06313_ sky130_fd_sc_hd__nor2_1
X_10963_ _03261_ _03264_ VGND VGND VPWR VPWR _03265_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12702_ _05174_ _05176_ VGND VGND VPWR VPWR _05177_ sky130_fd_sc_hd__nor2_1
XFILLER_0_57_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13682_ _06185_ _06236_ VGND VGND VPWR VPWR _06237_ sky130_fd_sc_hd__or2_2
X_10894_ _03187_ _03188_ VGND VGND VPWR VPWR _03189_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12794__B _02168_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12633_ _00392_ _02168_ _02723_ _00389_ VGND VGND VPWR VPWR _05101_ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_810 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12564_ _05013_ _05010_ VGND VGND VPWR VPWR _05025_ sky130_fd_sc_hd__nand2_1
XFILLER_0_109_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11515_ _03869_ _03870_ VGND VGND VPWR VPWR _03871_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire131 _01242_ VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__buf_2
XANTENNA__07400__C _03707_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12495_ _04037_ _03938_ VGND VGND VPWR VPWR _04949_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08215__D _00258_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11446_ _00262_ _03682_ _03678_ _00263_ VGND VGND VPWR VPWR _03796_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14165_ _06708_ _06735_ VGND VGND VPWR VPWR _06764_ sky130_fd_sc_hd__and2b_1
X_11377_ _03701_ _03719_ VGND VGND VPWR VPWR _03720_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13116_ _03456_ _03496_ _03625_ _03671_ VGND VGND VPWR VPWR _05633_ sky130_fd_sc_hd__o31a_1
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10328_ _05027_ _00373_ VGND VGND VPWR VPWR _02568_ sky130_fd_sc_hd__nand2_1
XANTENNA__07409__A _01197_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13489__B1 _01062_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14096_ _06645_ _06689_ _06690_ VGND VGND VPWR VPWR _06692_ sky130_fd_sc_hd__or3_4
XFILLER_0_147_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13047_ _05549_ _05556_ VGND VGND VPWR VPWR _05557_ sky130_fd_sc_hd__nand2_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10259_ _01833_ _02044_ _02052_ VGND VGND VPWR VPWR _02493_ sky130_fd_sc_hd__o21bai_1
XANTENNA__08904__A1 _00388_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08904__B2 _03004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10489__B _02743_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13949_ _06526_ _06529_ VGND VGND VPWR VPWR _06531_ sky130_fd_sc_hd__and2_1
XFILLER_0_76_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07470_ _01197_ _04367_ _04455_ _04510_ VGND VGND VPWR VPWR _04521_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09880__A2 _00416_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12216__A1 _01664_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12216__B2 _00607_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09140_ _01257_ _01202_ _01266_ VGND VGND VPWR VPWR _01267_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_29_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_284 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__10778__A1 _06937_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09071_ _00924_ _00927_ _01191_ VGND VGND VPWR VPWR _01192_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_127_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08022_ _00064_ _00065_ VGND VGND VPWR VPWR _00066_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09396__A1 _04169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_130_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09396__B2 _00431_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11767__C _01954_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09973_ _02175_ _02178_ VGND VGND VPWR VPWR _02179_ sky130_fd_sc_hd__xnor2_1
X_08924_ _00992_ _00839_ _01029_ VGND VGND VPWR VPWR _01031_ sky130_fd_sc_hd__and3_1
XFILLER_0_110_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08855_ _00773_ _00953_ VGND VGND VPWR VPWR _00955_ sky130_fd_sc_hd__or2_1
X_07806_ net148 net166 VGND VGND VPWR VPWR _06935_ sky130_fd_sc_hd__xnor2_2
XANTENNA__12598__C _01411_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08786_ _00707_ _00709_ VGND VGND VPWR VPWR _00881_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07737_ _00420_ net38 net37 net177 VGND VGND VPWR VPWR _06866_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07668_ _06658_ _06669_ VGND VGND VPWR VPWR _06680_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_1_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07204__D net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09407_ _01487_ _01490_ _01559_ VGND VGND VPWR VPWR _01560_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_94_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__13404__B1 _03687_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07882__A1 _00978_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07599_ _05901_ _05912_ VGND VGND VPWR VPWR _05923_ sky130_fd_sc_hd__nand2_1
XANTENNA__07882__B2 net149 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09338_ _01445_ _01446_ _01483_ VGND VGND VPWR VPWR _01484_ sky130_fd_sc_hd__or3_1
XFILLER_0_62_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09269_ _01407_ _01408_ VGND VGND VPWR VPWR _01409_ sky130_fd_sc_hd__or2_1
XFILLER_0_50_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11300_ _02785_ _03635_ VGND VGND VPWR VPWR _03636_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_90_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13707__A1 _02726_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12280_ _04711_ _04712_ VGND VGND VPWR VPWR _04713_ sky130_fd_sc_hd__or2b_1
XANTENNA__11958__B _02459_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11231_ _03556_ _03559_ VGND VGND VPWR VPWR _03560_ sky130_fd_sc_hd__or2_2
XFILLER_0_132_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11162_ _03470_ _03482_ _03483_ VGND VGND VPWR VPWR _03484_ sky130_fd_sc_hd__a21o_2
XANTENNA__09147__C _01272_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11396__D _02119_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10113_ _02321_ _02331_ VGND VGND VPWR VPWR _02332_ sky130_fd_sc_hd__xnor2_2
X_11093_ _03358_ _03407_ VGND VGND VPWR VPWR _03408_ sky130_fd_sc_hd__nor2_1
XANTENNA__09444__A _01586_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10044_ _01847_ _02255_ VGND VGND VPWR VPWR _02257_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13803_ _03414_ _03679_ _06369_ VGND VGND VPWR VPWR _06370_ sky130_fd_sc_hd__and3_1
X_11995_ _04392_ _04397_ _04396_ VGND VGND VPWR VPWR _04399_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_98_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output119_A net119 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12997__A2 _05494_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_836 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13734_ _00915_ _02725_ VGND VGND VPWR VPWR _06294_ sky130_fd_sc_hd__nand2_1
X_10946_ _03172_ _03187_ _03244_ VGND VGND VPWR VPWR _03247_ sky130_fd_sc_hd__o21a_1
XFILLER_0_42_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__09862__A2 _01188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_128_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13665_ _06216_ _06206_ VGND VGND VPWR VPWR _06218_ sky130_fd_sc_hd__or2b_1
X_10877_ _03093_ _03170_ VGND VGND VPWR VPWR _03171_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_66_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12616_ _05073_ _05080_ _05081_ VGND VGND VPWR VPWR _05083_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_109_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13596_ _06129_ _06141_ VGND VGND VPWR VPWR _06143_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12547_ _04978_ VGND VGND VPWR VPWR _05007_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12478_ _04915_ _04918_ VGND VGND VPWR VPWR _04931_ sky130_fd_sc_hd__or2_1
XFILLER_0_124_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14217_ _06803_ _02401_ VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__xnor2_2
XFILLER_0_112_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11429_ _03765_ _03767_ VGND VGND VPWR VPWR _03777_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14148_ _06729_ _06746_ VGND VGND VPWR VPWR _06747_ sky130_fd_sc_hd__or2b_1
XANTENNA__07139__A _00880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14079_ _06661_ _06672_ VGND VGND VPWR VPWR _06673_ sky130_fd_sc_hd__nand2_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08640_ _00565_ _00566_ _00569_ _00720_ VGND VGND VPWR VPWR _00721_ sky130_fd_sc_hd__or4_4
XANTENNA__09073__B _05731_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xrebuffer15 _00716_ VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__clkbuf_1
Xrebuffer26 net171 VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12211__C _01954_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer37 _03367_ VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__dlymetal6s2s_1
X_08571_ _06965_ _06966_ _00095_ _00151_ VGND VGND VPWR VPWR _00645_ sky130_fd_sc_hd__and4_1
XFILLER_0_49_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07522_ _03147_ net60 _00355_ _02960_ VGND VGND VPWR VPWR _05093_ sky130_fd_sc_hd__and4_1
XFILLER_0_76_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_735 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07453_ _04312_ _04323_ VGND VGND VPWR VPWR _04334_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_76_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13430__A_N _05424_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10666__C _02856_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07384_ _00431_ VGND VGND VPWR VPWR _03576_ sky130_fd_sc_hd__buf_4
XFILLER_0_17_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09123_ _01247_ VGND VGND VPWR VPWR _01248_ sky130_fd_sc_hd__buf_2
XFILLER_0_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09054_ _00557_ _01167_ _01172_ VGND VGND VPWR VPWR _01173_ sky130_fd_sc_hd__a21o_1
XFILLER_0_72_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08005_ _01044_ _03147_ _04367_ _04455_ VGND VGND VPWR VPWR _00049_ sky130_fd_sc_hd__nand4_1
XFILLER_0_13_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09956_ _02157_ _02159_ VGND VGND VPWR VPWR _02161_ sky130_fd_sc_hd__and2_1
X_08907_ _01010_ _01012_ VGND VGND VPWR VPWR _01013_ sky130_fd_sc_hd__or2_1
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09887_ _02082_ _02084_ VGND VGND VPWR VPWR _02085_ sky130_fd_sc_hd__or2_1
XANTENNA__12676__A1 _00381_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10687__B1 _02158_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08838_ _00751_ _00761_ VGND VGND VPWR VPWR _00937_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09414__D net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08769_ _00692_ _00860_ VGND VGND VPWR VPWR _00862_ sky130_fd_sc_hd__nor2_1
XFILLER_0_68_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10800_ _03074_ _03077_ VGND VGND VPWR VPWR _03086_ sky130_fd_sc_hd__or2_1
XFILLER_0_67_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11780_ _04161_ _04162_ VGND VGND VPWR VPWR _04163_ sky130_fd_sc_hd__nor2_1
XANTENNA__07304__B1 _00573_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10731_ _02989_ _03009_ VGND VGND VPWR VPWR _03010_ sky130_fd_sc_hd__or2_1
XFILLER_0_137_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__11034__A _00143_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13450_ _05969_ _02722_ VGND VGND VPWR VPWR _05982_ sky130_fd_sc_hd__nand2_1
XFILLER_0_137_256 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10662_ _02931_ _02928_ VGND VGND VPWR VPWR _02934_ sky130_fd_sc_hd__and2b_1
XFILLER_0_36_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12401_ _04834_ _04845_ VGND VGND VPWR VPWR _04846_ sky130_fd_sc_hd__nor2_1
XFILLER_0_51_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13381_ _05900_ _05906_ VGND VGND VPWR VPWR _05907_ sky130_fd_sc_hd__and2_1
XFILLER_0_118_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_788 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10593_ _02857_ VGND VGND VPWR VPWR _02858_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_63_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12332_ _04761_ _04769_ _04759_ VGND VGND VPWR VPWR _04770_ sky130_fd_sc_hd__o21a_1
XFILLER_0_105_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12263_ _04692_ _04693_ VGND VGND VPWR VPWR _04694_ sky130_fd_sc_hd__and2_1
XFILLER_0_121_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14002_ _06531_ _06523_ _06530_ VGND VGND VPWR VPWR _06589_ sky130_fd_sc_hd__or3_1
X_11214_ _03539_ _03540_ VGND VGND VPWR VPWR _03541_ sky130_fd_sc_hd__and2_1
X_12194_ _04617_ _04613_ VGND VGND VPWR VPWR _04618_ sky130_fd_sc_hd__or2_1
Xoutput73 net73 VGND VGND VPWR VPWR prod[17] sky130_fd_sc_hd__clkbuf_4
X_11145_ _03461_ _03462_ _03464_ VGND VGND VPWR VPWR _03465_ sky130_fd_sc_hd__a21o_1
Xoutput84 net84 VGND VGND VPWR VPWR prod[27] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput95 net95 VGND VGND VPWR VPWR prod[37] sky130_fd_sc_hd__buf_2
X_11076_ _03330_ _03326_ _03328_ VGND VGND VPWR VPWR _03390_ sky130_fd_sc_hd__nor3_1
XANTENNA__12312__B _00607_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10027_ _01916_ _01939_ _02238_ VGND VGND VPWR VPWR _02239_ sky130_fd_sc_hd__o21a_1
XFILLER_0_144_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11978_ _04377_ _04379_ VGND VGND VPWR VPWR _04381_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10929_ _03212_ _03227_ VGND VGND VPWR VPWR _03228_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13717_ _06270_ _06275_ VGND VGND VPWR VPWR _06276_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_711 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_839 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07141__B _00901_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13648_ _06196_ _06199_ VGND VGND VPWR VPWR _06200_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13579_ _06122_ _06123_ VGND VGND VPWR VPWR _06124_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09349__A _05192_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09068__B _01188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09810_ _01998_ _02000_ VGND VGND VPWR VPWR _02001_ sky130_fd_sc_hd__nor2_1
XANTENNA__12503__A _00378_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__08700__B _00779_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09741_ _04268_ net50 VGND VGND VPWR VPWR _01925_ sky130_fd_sc_hd__nand2_1
X_09672_ _01847_ _01848_ VGND VGND VPWR VPWR _01849_ sky130_fd_sc_hd__nor2_1
XANTENNA__08371__A2_N net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08623_ _00513_ _00701_ VGND VGND VPWR VPWR _00702_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_11_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08554_ _00624_ _00625_ VGND VGND VPWR VPWR _00626_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10677__B _01411_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07332__A _02993_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07505_ _04895_ VGND VGND VPWR VPWR _04906_ sky130_fd_sc_hd__clkbuf_4
X_08485_ _00465_ _00549_ _00548_ VGND VGND VPWR VPWR _00551_ sky130_fd_sc_hd__o21a_1
XFILLER_0_65_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07436_ _04092_ _04136_ VGND VGND VPWR VPWR _04147_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09039__B1 _01155_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_119_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12892__B _02459_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07367_ _03246_ _03378_ VGND VGND VPWR VPWR _03389_ sky130_fd_sc_hd__xor2_1
XFILLER_0_33_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11397__A1 _00112_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09106_ _00530_ _00391_ _01228_ VGND VGND VPWR VPWR _01231_ sky130_fd_sc_hd__a21o_1
XANTENNA__11397__B2 _00268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13500__C _01415_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07298_ net169 _02620_ VGND VGND VPWR VPWR _02631_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09037_ _00544_ VGND VGND VPWR VPWR _01155_ sky130_fd_sc_hd__buf_4
XFILLER_0_130_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__07507__A _04873_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09939_ _02111_ _02141_ VGND VGND VPWR VPWR _02142_ sky130_fd_sc_hd__nor2_1
X_12950_ _05024_ _05026_ VGND VGND VPWR VPWR _05450_ sky130_fd_sc_hd__nor2_2
X_11901_ _02280_ _03678_ _04295_ VGND VGND VPWR VPWR _04296_ sky130_fd_sc_hd__and3_1
XTAP_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12881_ _05372_ _05373_ VGND VGND VPWR VPWR _05374_ sky130_fd_sc_hd__xnor2_1
XTAP_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11872__A2 _01780_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09441__B _02018_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11832_ _04186_ _02677_ _04187_ VGND VGND VPWR VPWR _04220_ sky130_fd_sc_hd__a21oi_1
XTAP_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08338__A _00390_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07242__A _02007_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07828__A1 _00880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11763_ _00138_ _01953_ _02134_ _02018_ VGND VGND VPWR VPWR _04144_ sky130_fd_sc_hd__a22o_1
XTAP_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13502_ _06037_ _06038_ VGND VGND VPWR VPWR _06039_ sky130_fd_sc_hd__nor2_1
X_10714_ _02939_ _02948_ _02989_ _02937_ VGND VGND VPWR VPWR _02991_ sky130_fd_sc_hd__o31ai_2
XTAP_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11694_ _04062_ _04067_ VGND VGND VPWR VPWR _04068_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13433_ _05422_ _05963_ VGND VGND VPWR VPWR _05964_ sky130_fd_sc_hd__and2_1
XANTENNA__07896__B _03499_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10645_ _02913_ _02914_ VGND VGND VPWR VPWR _02915_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__12585__B1 _02304_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13364_ _01289_ _02759_ _02721_ _02008_ VGND VGND VPWR VPWR _05888_ sky130_fd_sc_hd__a22o_1
Xrebuffer6 _02576_ VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_63_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10576_ _02829_ _02826_ VGND VGND VPWR VPWR _02840_ sky130_fd_sc_hd__and2b_1
XFILLER_0_90_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12315_ _00608_ _01601_ _04737_ _04738_ VGND VGND VPWR VPWR _04751_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_133_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13295_ _05696_ _05711_ VGND VGND VPWR VPWR _05817_ sky130_fd_sc_hd__and2b_1
XFILLER_0_23_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12246_ _04037_ _00783_ _01178_ _01248_ VGND VGND VPWR VPWR _04676_ sky130_fd_sc_hd__and4_1
XFILLER_0_139_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12177_ _04024_ net186 _04597_ _04599_ VGND VGND VPWR VPWR _04600_ sky130_fd_sc_hd__o211a_4
X_11128_ _03386_ _03402_ _03441_ _03445_ _03446_ VGND VGND VPWR VPWR _03447_ sky130_fd_sc_hd__a41o_1
XANTENNA__07417__A net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11059_ _03369_ _03370_ VGND VGND VPWR VPWR _03371_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07152__A net1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08270_ _00148_ _00315_ VGND VGND VPWR VPWR _00316_ sky130_fd_sc_hd__nand2_1
XFILLER_0_144_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07221_ _01766_ _01777_ VGND VGND VPWR VPWR _01788_ sky130_fd_sc_hd__nor2_4
XFILLER_0_104_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_861 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_703 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07152_ net1 net62 net12 net61 VGND VGND VPWR VPWR _01033_ sky130_fd_sc_hd__and4_1
XFILLER_0_82_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_739 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10960__B _00310_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11000__B1 _00959_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07985_ _07020_ _07027_ VGND VGND VPWR VPWR _00029_ sky130_fd_sc_hd__and2_1
X_09724_ _01904_ _01905_ VGND VGND VPWR VPWR _01906_ sky130_fd_sc_hd__or2_1
X_09655_ _01626_ _01561_ _01560_ VGND VGND VPWR VPWR _01831_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_97_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__10688__A _00366_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08606_ _00681_ _00682_ VGND VGND VPWR VPWR _00684_ sky130_fd_sc_hd__nor2_1
XFILLER_0_145_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09586_ _01355_ _01486_ VGND VGND VPWR VPWR _01756_ sky130_fd_sc_hd__nor2_2
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08537_ _00607_ VGND VGND VPWR VPWR _00608_ sky130_fd_sc_hd__buf_4
XFILLER_0_49_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__10200__B _02427_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_198 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08468_ _02993_ _06873_ _06875_ _05203_ VGND VGND VPWR VPWR _00533_ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07419_ _03927_ _03949_ VGND VGND VPWR VPWR _03960_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_179 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08399_ net45 VGND VGND VPWR VPWR _00457_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_80_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10430_ _02466_ _02679_ VGND VGND VPWR VPWR _02680_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_864 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10361_ _02602_ _02603_ VGND VGND VPWR VPWR _02604_ sky130_fd_sc_hd__xor2_1
XFILLER_0_115_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12100_ _04503_ _04514_ VGND VGND VPWR VPWR _04515_ sky130_fd_sc_hd__xnor2_2
XANTENNA__11790__A1 _01295_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11790__B2 _01306_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13080_ _05545_ _05592_ _05543_ VGND VGND VPWR VPWR _05593_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_103_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10292_ _02526_ _02527_ VGND VGND VPWR VPWR _02528_ sky130_fd_sc_hd__xor2_1
XFILLER_0_103_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12031_ _04428_ _04438_ VGND VGND VPWR VPWR _04439_ sky130_fd_sc_hd__and2b_1
XANTENNA__08538__A2 _00458_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__10345__A2 _02377_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13819__B1 _03686_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13982_ _06553_ _06566_ VGND VGND VPWR VPWR _06567_ sky130_fd_sc_hd__nor2_1
X_12933_ _03585_ _03588_ _03590_ VGND VGND VPWR VPWR _05431_ sky130_fd_sc_hd__and3_2
XFILLER_0_87_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13405__C _01955_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__08068__A _07010_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12864_ _05292_ _05354_ VGND VGND VPWR VPWR _05355_ sky130_fd_sc_hd__nand2_1
XTAP_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_817 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11815_ _04199_ _04200_ VGND VGND VPWR VPWR _04201_ sky130_fd_sc_hd__nor2_1
XFILLER_0_139_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output101_A net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12795_ _05277_ _05278_ VGND VGND VPWR VPWR _05279_ sky130_fd_sc_hd__xor2_1
XTAP_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11746_ _00543_ _01188_ VGND VGND VPWR VPWR _04126_ sky130_fd_sc_hd__nand2_1
XTAP_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12270__A2 _01181_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11677_ _07010_ _03773_ _01260_ _00268_ VGND VGND VPWR VPWR _04050_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08226__A1 _02116_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10628_ _02813_ _02841_ VGND VGND VPWR VPWR _02897_ sky130_fd_sc_hd__nor2_1
X_13416_ _05853_ _05943_ _05944_ VGND VGND VPWR VPWR _05946_ sky130_fd_sc_hd__and3_1
XFILLER_0_24_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08226__B2 _02149_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13347_ _05342_ _05345_ _05343_ VGND VGND VPWR VPWR _05870_ sky130_fd_sc_hd__o21ba_1
X_10559_ _02819_ _02820_ VGND VGND VPWR VPWR _02821_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_11_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10584__A2 _02306_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13278_ _05472_ _05732_ VGND VGND VPWR VPWR _05801_ sky130_fd_sc_hd__and2_1
XFILLER_0_11_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12229_ _01518_ _03750_ VGND VGND VPWR VPWR _04657_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_794 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07737__B1 net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07147__A net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07770_ _05412_ _06897_ _06898_ VGND VGND VPWR VPWR _06899_ sky130_fd_sc_hd__o21bai_2
XANTENNA__09362__A _01350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09440_ _01573_ _01595_ VGND VGND VPWR VPWR _01596_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_91_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09371_ _06483_ _01517_ _01519_ VGND VGND VPWR VPWR _01520_ sky130_fd_sc_hd__and3_2
X_08322_ _04015_ VGND VGND VPWR VPWR _00373_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08253_ _00163_ _00162_ VGND VGND VPWR VPWR _00297_ sky130_fd_sc_hd__and2b_1
XFILLER_0_6_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07967__D net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07204_ _00420_ _00978_ _01208_ net44 VGND VGND VPWR VPWR _01602_ sky130_fd_sc_hd__and4_1
XFILLER_0_144_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08184_ _00221_ _00227_ VGND VGND VPWR VPWR _00228_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_27_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09965__A1 _02051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07135_ net153 _00836_ VGND VGND VPWR VPWR _00847_ sky130_fd_sc_hd__or2b_1
XANTENNA__09965__B2 _00453_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10971__A _00142_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__09537__A _05192_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07968_ _00010_ _00011_ VGND VGND VPWR VPWR _00012_ sky130_fd_sc_hd__nand2_1
XANTENNA__09272__A _01411_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09707_ _01885_ _01887_ VGND VGND VPWR VPWR _01888_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07899_ _07020_ _07027_ VGND VGND VPWR VPWR _07028_ sky130_fd_sc_hd__xor2_1
XFILLER_0_97_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09638_ _01811_ _01812_ VGND VGND VPWR VPWR _01813_ sky130_fd_sc_hd__xor2_1
XFILLER_0_78_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09569_ _01735_ _01736_ VGND VGND VPWR VPWR _01737_ sky130_fd_sc_hd__and2_1
XFILLER_0_84_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11600_ _03827_ _03829_ VGND VGND VPWR VPWR _03965_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12580_ _03740_ _00742_ _02849_ _02304_ VGND VGND VPWR VPWR _05043_ sky130_fd_sc_hd__and4_1
XFILLER_0_136_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11531_ _03877_ _03888_ VGND VGND VPWR VPWR _03889_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_65_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__11042__A _00158_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11462_ _00121_ net21 _02133_ _03521_ VGND VGND VPWR VPWR _03813_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10156__B1_N _02235_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13201_ _05457_ _05469_ VGND VGND VPWR VPWR _05726_ sky130_fd_sc_hd__and2_1
X_10413_ _02454_ _02659_ VGND VGND VPWR VPWR _02661_ sky130_fd_sc_hd__and2_1
X_14181_ _06761_ _06762_ _06779_ _06780_ VGND VGND VPWR VPWR _06781_ sky130_fd_sc_hd__a211o_1
X_11393_ _00113_ _01179_ _01249_ _00114_ VGND VGND VPWR VPWR _03737_ sky130_fd_sc_hd__a22oi_1
XANTENNA__11763__A1 _00138_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13132_ _05609_ _05615_ _05617_ _04031_ VGND VGND VPWR VPWR _05650_ sky130_fd_sc_hd__or4_1
XFILLER_0_103_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11763__B2 _02018_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10344_ _02334_ _02345_ VGND VGND VPWR VPWR _02585_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_571 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_284 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13063_ _05572_ _05568_ _05570_ VGND VGND VPWR VPWR _05574_ sky130_fd_sc_hd__and3_1
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10275_ net57 _02507_ _02508_ VGND VGND VPWR VPWR _02509_ sky130_fd_sc_hd__a21bo_1
XANTENNA__12304__C _00608_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12014_ _04418_ _04408_ VGND VGND VPWR VPWR _04420_ sky130_fd_sc_hd__and2b_1
XANTENNA__07195__A1 _00420_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10105__B _05742_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07195__B2 _00978_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13965_ _06349_ _05897_ _06350_ VGND VGND VPWR VPWR _06548_ sky130_fd_sc_hd__nand3_1
XANTENNA__07414__B _03894_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12916_ _05304_ _05410_ _05409_ VGND VGND VPWR VPWR _05413_ sky130_fd_sc_hd__a21o_1
XANTENNA__12491__A2 _03696_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13896_ _05363_ _05405_ _05941_ VGND VGND VPWR VPWR _06473_ sky130_fd_sc_hd__or3_1
XTAP_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12847_ _05334_ _05336_ VGND VGND VPWR VPWR _05337_ sky130_fd_sc_hd__and2_1
XTAP_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12778_ _04775_ _05037_ VGND VGND VPWR VPWR _05261_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__11673__A2_N _03938_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__07430__A _01284_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__13151__B _05670_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11729_ _04055_ _02608_ _04056_ VGND VGND VPWR VPWR _04107_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11203__B1 _03503_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_142_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09357__A _01504_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08940_ _00984_ _01048_ VGND VGND VPWR VPWR _01049_ sky130_fd_sc_hd__xor2_2
XANTENNA__08723__A2_N _00144_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08871_ _00787_ _00788_ VGND VGND VPWR VPWR _00973_ sky130_fd_sc_hd__nand2_1
X_07822_ _06949_ _06950_ VGND VGND VPWR VPWR _06951_ sky130_fd_sc_hd__or2_1
XANTENNA__13607__A _01061_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_07753_ _06864_ _06881_ VGND VGND VPWR VPWR _06882_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11772__D net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12230__B _03748_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07684_ net12 net35 net34 net149 VGND VGND VPWR VPWR _06813_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09423_ _06417_ _00745_ _01575_ _01263_ VGND VGND VPWR VPWR _01577_ sky130_fd_sc_hd__a31o_1
XANTENNA__11690__B1 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09354_ _01380_ _01393_ VGND VGND VPWR VPWR _01501_ sky130_fd_sc_hd__nand2_1
XANTENNA__08436__A _05478_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__12234__A2 _01178_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13699__D _02720_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08305_ _04158_ _00353_ VGND VGND VPWR VPWR _00354_ sky130_fd_sc_hd__nand2_2
XANTENNA__07340__A _02007_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__11442__B1 _02459_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09285_ _01359_ _01425_ VGND VGND VPWR VPWR _01426_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_47_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_80 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08236_ _00108_ _00279_ VGND VGND VPWR VPWR _00280_ sky130_fd_sc_hd__nor2_1
XFILLER_0_145_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08167_ net167 _06076_ VGND VGND VPWR VPWR _00211_ sky130_fd_sc_hd__or2b_1
XANTENNA__10548__A2 _02725_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07118_ net44 VGND VGND VPWR VPWR _00661_ sky130_fd_sc_hd__buf_6
X_08098_ _05027_ VGND VGND VPWR VPWR _00142_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_30_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10060_ _01837_ _02045_ VGND VGND VPWR VPWR _02275_ sky130_fd_sc_hd__and2_1
XANTENNA__07218__C _01744_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10579__C _02306_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10962_ _03262_ _03263_ VGND VGND VPWR VPWR _03264_ sky130_fd_sc_hd__nor2_1
X_13750_ _06309_ _06310_ VGND VGND VPWR VPWR _06312_ sky130_fd_sc_hd__and2_1
XFILLER_0_98_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12701_ _05078_ _05175_ VGND VGND VPWR VPWR _05176_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13681_ _06189_ _06235_ VGND VGND VPWR VPWR _06236_ sky130_fd_sc_hd__nor2_1
X_10893_ _03174_ _03186_ VGND VGND VPWR VPWR _03188_ sky130_fd_sc_hd__and2_1
XANTENNA__13252__A _05546_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12632_ _00389_ _00392_ _02723_ VGND VGND VPWR VPWR _05100_ sky130_fd_sc_hd__and3_1
XFILLER_0_38_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_822 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__07250__A _00628_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12563_ _05021_ _05023_ VGND VGND VPWR VPWR _05024_ sky130_fd_sc_hd__nand2_2
XFILLER_0_93_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_628 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11514_ _03865_ _03867_ VGND VGND VPWR VPWR _03870_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12494_ _04936_ _04935_ VGND VGND VPWR VPWR _04948_ sky130_fd_sc_hd__and2b_1
XFILLER_0_108_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07400__D _03740_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14233_ _06811_ _06807_ VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__xnor2_2
X_11445_ _00262_ _00263_ _03682_ _03679_ VGND VGND VPWR VPWR _03794_ sky130_fd_sc_hd__nand4_1
XFILLER_0_123_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14164_ _06761_ _06762_ VGND VGND VPWR VPWR _06763_ sky130_fd_sc_hd__xor2_1
X_11376_ _03695_ _03698_ _03700_ _03692_ VGND VGND VPWR VPWR _03719_ sky130_fd_sc_hd__o22a_1
XFILLER_0_22_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10327_ _00613_ _02564_ _02566_ VGND VGND VPWR VPWR _02567_ sky130_fd_sc_hd__a21bo_1
X_13115_ _05628_ _05630_ VGND VGND VPWR VPWR _05631_ sky130_fd_sc_hd__xor2_2
X_14095_ _06610_ _06628_ VGND VGND VPWR VPWR _06690_ sky130_fd_sc_hd__or2_1
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13046_ _05551_ _05554_ VGND VGND VPWR VPWR _05556_ sky130_fd_sc_hd__nor2_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10258_ _02045_ _02274_ VGND VGND VPWR VPWR _02492_ sky130_fd_sc_hd__and2_2
XANTENNA__08904__A2 _00112_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10189_ _02414_ _00734_ _00486_ _02411_ VGND VGND VPWR VPWR _02416_ sky130_fd_sc_hd__and4b_1
XANTENNA__07425__A _04015_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13948_ _06526_ _06529_ VGND VGND VPWR VPWR _06530_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09640__A _00311_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13879_ _05913_ _05927_ VGND VGND VPWR VPWR _06454_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12216__A2 _01180_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__07160__A net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10778__A2 _02169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09070_ _00925_ _00926_ VGND VGND VPWR VPWR _01191_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08021_ _00058_ _00063_ VGND VGND VPWR VPWR _00065_ sky130_fd_sc_hd__and2_1
XFILLER_0_72_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__09396__A2 net50 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_142_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__11767__D _02135_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_122_390 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09972_ _02176_ _02177_ VGND VGND VPWR VPWR _02178_ sky130_fd_sc_hd__nor2_1
XFILLER_0_110_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08923_ _00992_ _00839_ _01029_ VGND VGND VPWR VPWR _01030_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07159__A1 _00880_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08854_ _00773_ _00953_ VGND VGND VPWR VPWR _00954_ sky130_fd_sc_hd__nand2_1
XANTENNA__07335__A _01470_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07805_ _05302_ _05368_ _05390_ _06933_ VGND VGND VPWR VPWR _06934_ sky130_fd_sc_hd__o31ai_2
XANTENNA__12598__D _02849_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08785_ _00553_ _00556_ _00710_ VGND VGND VPWR VPWR _00879_ sky130_fd_sc_hd__or3_1
XFILLER_0_137_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07736_ _00420_ net177 net38 net37 VGND VGND VPWR VPWR _06865_ sky130_fd_sc_hd__and4_1
XANTENNA__12895__B _02673_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07667_ _06263_ _06549_ _06582_ VGND VGND VPWR VPWR _06669_ sky130_fd_sc_hd__a21o_1
XANTENNA__11663__B1 _00574_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09406_ _01423_ _01557_ VGND VGND VPWR VPWR _01559_ sky130_fd_sc_hd__xor2_1
XFILLER_0_1_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__13404__A1 _03414_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07598_ _05857_ _05890_ VGND VGND VPWR VPWR _05912_ sky130_fd_sc_hd__or2_1
XANTENNA__07882__A2 _07010_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__13404__B2 _04714_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10218__A1 _05731_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10218__B2 _01000_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09337_ _01479_ _01482_ VGND VGND VPWR VPWR _01483_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13800__A _02187_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09268_ _01064_ _01105_ _01406_ VGND VGND VPWR VPWR _01408_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_106_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08219_ _06966_ VGND VGND VPWR VPWR _00263_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_62_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09199_ _01137_ _01140_ VGND VGND VPWR VPWR _01332_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__12416__A _00378_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11230_ _03557_ _03558_ VGND VGND VPWR VPWR _03559_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__08595__B1 _00670_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11161_ _03471_ _03481_ VGND VGND VPWR VPWR _03483_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__09147__D _01211_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10112_ _02329_ _02330_ VGND VGND VPWR VPWR _02331_ sky130_fd_sc_hd__nor2_1
X_11092_ _02574_ _03357_ VGND VGND VPWR VPWR _03407_ sky130_fd_sc_hd__and2_1
X_10043_ _01847_ _02255_ VGND VGND VPWR VPWR _02256_ sky130_fd_sc_hd__and2_1
XANTENNA__07245__A _00989_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13802_ _06366_ _06368_ VGND VGND VPWR VPWR _06369_ sky130_fd_sc_hd__nor2_1
X_11994_ _04392_ _04396_ _04397_ VGND VGND VPWR VPWR _04398_ sky130_fd_sc_hd__or3_4
XFILLER_0_98_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13733_ _05855_ _05859_ VGND VGND VPWR VPWR _06293_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10945_ _03244_ _03172_ VGND VGND VPWR VPWR _03245_ sky130_fd_sc_hd__or2_1
XFILLER_0_86_848 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13664_ _06206_ _06216_ VGND VGND VPWR VPWR _06217_ sky130_fd_sc_hd__or2b_1
XFILLER_0_128_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10876_ _03099_ _03098_ VGND VGND VPWR VPWR _03170_ sky130_fd_sc_hd__or2b_1
XANTENNA__11214__B _03540_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12615_ _05065_ _05070_ _05072_ VGND VGND VPWR VPWR _05081_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_66_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13595_ _06127_ _06128_ _06126_ VGND VGND VPWR VPWR _06141_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_26_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__13710__A _02759_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_124_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12546_ _00393_ _00459_ _01400_ _00390_ VGND VGND VPWR VPWR _05006_ sky130_fd_sc_hd__a22o_1
XFILLER_0_124_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12477_ _04714_ _02008_ VGND VGND VPWR VPWR _04930_ sky130_fd_sc_hd__and2_1
XANTENNA__12326__A _00460_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__11868__C _00003_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output93_A net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14216_ _02412_ _02248_ VGND VGND VPWR VPWR _06803_ sky130_fd_sc_hd__or2b_1
X_11428_ _03774_ _03775_ VGND VGND VPWR VPWR _03776_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14147_ _06743_ _06745_ VGND VGND VPWR VPWR _06746_ sky130_fd_sc_hd__nand2_1
X_11359_ _01155_ _03699_ _03691_ VGND VGND VPWR VPWR _03700_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14078_ _06666_ _06671_ VGND VGND VPWR VPWR _06672_ sky130_fd_sc_hd__xnor2_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13029_ _02589_ _04604_ _03551_ VGND VGND VPWR VPWR _05537_ sky130_fd_sc_hd__o21ai_2
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09073__C _03718_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xrebuffer16 net163 VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__clkbuf_1
X_08570_ _06965_ _00293_ _00151_ _00263_ VGND VGND VPWR VPWR _00644_ sky130_fd_sc_hd__a22oi_1
Xrebuffer27 _07047_ VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__12211__D _02135_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xrebuffer38 _02740_ VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_77_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__09370__A _06461_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07521_ _05060_ _05071_ VGND VGND VPWR VPWR _05082_ sky130_fd_sc_hd__and2_1
XFILLER_0_88_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07452_ _04158_ _04301_ VGND VGND VPWR VPWR _04323_ sky130_fd_sc_hd__nand2_1
XANTENNA__11405__A _02119_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_147_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__10666__D _02858_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07383_ _00453_ _03554_ _00519_ _02051_ VGND VGND VPWR VPWR _03565_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_44_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09122_ _01246_ VGND VGND VPWR VPWR _01247_ sky130_fd_sc_hd__buf_2
XFILLER_0_17_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09053_ _01170_ _01171_ VGND VGND VPWR VPWR _01172_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08004_ _01044_ _04367_ net3 _03147_ VGND VGND VPWR VPWR _00048_ sky130_fd_sc_hd__a22o_1
XFILLER_0_25_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_686 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09955_ _04081_ _01339_ _02158_ _02156_ VGND VGND VPWR VPWR _02159_ sky130_fd_sc_hd__nand4_2
X_08906_ _00003_ _00095_ _01008_ _01009_ VGND VGND VPWR VPWR _01012_ sky130_fd_sc_hd__o2bb2a_1
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09886_ _02058_ _02081_ VGND VGND VPWR VPWR _02084_ sky130_fd_sc_hd__and2_1
XANTENNA__12676__A2 _01958_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10687__A1 _02982_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__10687__B2 _00366_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08837_ _00913_ _00935_ VGND VGND VPWR VPWR _00936_ sky130_fd_sc_hd__xor2_4
X_08768_ _00692_ _00860_ VGND VGND VPWR VPWR _00861_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07719_ _06833_ _06839_ _06840_ VGND VGND VPWR VPWR _06848_ sky130_fd_sc_hd__o21a_1
X_08699_ _01383_ _00784_ VGND VGND VPWR VPWR _00785_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__07304__B2 net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10730_ _02988_ _02959_ _02987_ VGND VGND VPWR VPWR _03009_ sky130_fd_sc_hd__nor3_1
XFILLER_0_67_358 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10661_ _02920_ _02932_ VGND VGND VPWR VPWR _02933_ sky130_fd_sc_hd__xor2_4
XANTENNA__11034__B _01518_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_419 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12400_ _04832_ _04833_ _04831_ VGND VGND VPWR VPWR _04845_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_35_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13380_ _05902_ _05905_ VGND VGND VPWR VPWR _05906_ sky130_fd_sc_hd__xor2_1
X_10592_ _02305_ VGND VGND VPWR VPWR _02857_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_118_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10611__A1 _00310_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12331_ _04767_ _04768_ VGND VGND VPWR VPWR _04769_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12262_ _04681_ _04683_ VGND VGND VPWR VPWR _04693_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_121_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14001_ _06531_ _06530_ _06523_ VGND VGND VPWR VPWR _06588_ sky130_fd_sc_hd__o21ai_1
X_11213_ _03434_ _03436_ VGND VGND VPWR VPWR _03540_ sky130_fd_sc_hd__xor2_2
XFILLER_0_121_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__13561__B1 _02736_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12193_ _04614_ _04608_ _04616_ VGND VGND VPWR VPWR _04617_ sky130_fd_sc_hd__o21ba_1
XANTENNA__10375__B1 _00571_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11144_ _03045_ _03463_ VGND VGND VPWR VPWR _03464_ sky130_fd_sc_hd__nor2_2
Xoutput74 net74 VGND VGND VPWR VPWR prod[18] sky130_fd_sc_hd__clkbuf_4
Xoutput85 net85 VGND VGND VPWR VPWR prod[28] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_128_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput96 net96 VGND VGND VPWR VPWR prod[38] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11075_ _03373_ _03387_ VGND VGND VPWR VPWR _03388_ sky130_fd_sc_hd__xor2_1
XANTENNA__12312__C _01664_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10026_ _01916_ _01939_ _01889_ VGND VGND VPWR VPWR _02238_ sky130_fd_sc_hd__a21o_1
XFILLER_0_53_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11977_ _04377_ _04379_ VGND VGND VPWR VPWR _04380_ sky130_fd_sc_hd__nor2_1
XFILLER_0_129_703 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13716_ _06272_ _06273_ VGND VGND VPWR VPWR _06275_ sky130_fd_sc_hd__nor2_1
X_10928_ _03209_ _03211_ VGND VGND VPWR VPWR _03227_ sky130_fd_sc_hd__or2_1
XFILLER_0_129_747 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__10850__A1 _05566_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13647_ _06198_ _06016_ VGND VGND VPWR VPWR _06199_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10859_ _03268_ _01410_ VGND VGND VPWR VPWR _03151_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__08534__A net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13578_ _01250_ _02858_ _06121_ VGND VGND VPWR VPWR _06123_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_26_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__09349__B net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12529_ _04984_ _04986_ VGND VGND VPWR VPWR _04987_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__12503__B _00741_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09740_ _01922_ _01923_ VGND VGND VPWR VPWR _01924_ sky130_fd_sc_hd__nor2_1
.ends

