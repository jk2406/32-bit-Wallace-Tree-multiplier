// This is the unpowered netlist.
module wallacetree32x32 (a,
    b,
    prod);
 input [31:0] a;
 input [31:0] b;
 output [63:0] prod;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__diode_2 ANTENNA__07085__A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__07086__A (.DIODE(_00300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07087__A (.DIODE(_00311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07088__A (.DIODE(_00322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07089__A (.DIODE(_00333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07090__A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__07091__A (.DIODE(_00355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07092__A (.DIODE(_00366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07093__A (.DIODE(_00377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07094__A (.DIODE(_00388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07095__A (.DIODE(_00399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07096__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07097__A (.DIODE(_00420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07098__A (.DIODE(_00431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07099__A (.DIODE(_00442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07100__A (.DIODE(_00453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07101__A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__07102__A (.DIODE(_00475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07103__A (.DIODE(_00486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07104__A (.DIODE(_00497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07105__A (.DIODE(_00508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07106__A (.DIODE(_00519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07107__A (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__07108__A (.DIODE(_00541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07108__B (.DIODE(_00300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07109__A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__07110__A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__07111__A (.DIODE(_00563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07111__B (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__07111__C (.DIODE(_00573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07111__D (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__07112__A1 (.DIODE(_00563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07112__A2 (.DIODE(_00573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07112__B1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__07112__B2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__07115__A (.DIODE(_00563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07116__A (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__07117__A (.DIODE(_00639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07118__A (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__07119__A (.DIODE(_00661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07120__A (.DIODE(_00628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07120__B (.DIODE(_00650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07120__C (.DIODE(_00672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07120__D (.DIODE(_00300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07122__A (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__07123__A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__07124__A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__07124__C (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__07125__A1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__07125__B1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__07125__B2 (.DIODE(_00573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07127__A (.DIODE(_00541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07127__B (.DIODE(_00661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07129__A1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__07129__A2 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__07130__A (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__07130__B (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__07137__A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__07138__A (.DIODE(_00869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07139__A (.DIODE(_00880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07140__A (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__07141__A (.DIODE(_00891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07141__B (.DIODE(_00901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07142__A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__07143__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07143__C (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__07143__D (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__07144__A1 (.DIODE(_00420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07144__A2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__07144__B1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__07147__A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__07148__A (.DIODE(_00978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07149__A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__07150__A (.DIODE(_00442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07150__B (.DIODE(_00989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07150__C (.DIODE(_01000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07150__D (.DIODE(_00901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07152__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07152__B (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__07152__C (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__07152__D (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__07153__A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__07154__A1 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07154__A2 (.DIODE(_01044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07154__B2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__07156__A (.DIODE(_00869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07157__A (.DIODE(_01076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07157__B (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__07159__A1 (.DIODE(_00880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07159__A2 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__07160__A (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__07161__A (.DIODE(_01120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07161__B (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__07167__A (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__07169__A (.DIODE(_00880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07169__B (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__07169__C (.DIODE(_01197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07169__D (.DIODE(_01208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07170__A (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__07171__A1 (.DIODE(_00978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07171__B1 (.DIODE(_01208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07171__B2 (.DIODE(_00869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07172__B (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__07172__D (.DIODE(_00573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07173__A1 (.DIODE(_01230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07173__A2 (.DIODE(_00672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07175__A (.DIODE(_01076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07176__A (.DIODE(_01197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07177__A (.DIODE(_01208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07178__A1 (.DIODE(_01284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07178__A2 (.DIODE(_01295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07178__B1 (.DIODE(_01306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07178__B2 (.DIODE(_01230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07180__A (.DIODE(_01230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07181__A (.DIODE(_01339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07182__A (.DIODE(_01295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07183__A (.DIODE(_00891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07184__A (.DIODE(_01372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07185__A (.DIODE(_01208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07187__A (.DIODE(_01383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07187__B (.DIODE(_01405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07188__A (.DIODE(_01350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07188__B (.DIODE(_01361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07192__A (.DIODE(_00661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07193__A (.DIODE(_01120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07193__B (.DIODE(_01470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07195__A1 (.DIODE(_00420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07195__A2 (.DIODE(_01197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07195__B1 (.DIODE(_01208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07195__B2 (.DIODE(_00978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07196__A (.DIODE(_00420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07196__B (.DIODE(_00978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07196__D (.DIODE(_01208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07197__A1 (.DIODE(_01284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07197__A2 (.DIODE(_00672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07202__A (.DIODE(_01230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07202__B (.DIODE(_00300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07203__A1 (.DIODE(_00420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07203__A2 (.DIODE(_01208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07203__B1 (.DIODE(_00661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07203__B2 (.DIODE(_00978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07204__A (.DIODE(_00420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07204__B (.DIODE(_00978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07204__C (.DIODE(_01208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07204__D (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__07205__A1 (.DIODE(_01076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07205__A2 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__07208__A (.DIODE(_00891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07208__B (.DIODE(_00672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07215__A (.DIODE(_01284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07215__B (.DIODE(_00300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07217__A (.DIODE(_00672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07218__A (.DIODE(_00442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07218__B (.DIODE(_00989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07218__C (.DIODE(_01744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07218__D (.DIODE(_00311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07240__A (.DIODE(_01000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07241__A (.DIODE(_01996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07242__A (.DIODE(_02007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07243__A (.DIODE(_00901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07244__A (.DIODE(_02029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07245__A (.DIODE(_00989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07246__A1 (.DIODE(_00442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07246__A2 (.DIODE(_02018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07246__B1 (.DIODE(_02040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07246__B2 (.DIODE(_02051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07250__A (.DIODE(_00628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07251__A (.DIODE(_02105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07252__A (.DIODE(_00672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07253__A (.DIODE(_02127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07254__A (.DIODE(_00650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07255__A (.DIODE(_02149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07257__A1 (.DIODE(_02116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07257__A2 (.DIODE(_02138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07257__B1 (.DIODE(_00333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07257__B2 (.DIODE(_02171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07264__A (.DIODE(_02116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07265__A (.DIODE(_02259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07265__B (.DIODE(_00333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07266__A (.DIODE(_02040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07270__A (.DIODE(_00453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07270__B (.DIODE(_02280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07271__A (.DIODE(_02280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07272__A1 (.DIODE(_00453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07272__A2 (.DIODE(_02335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07282__A (.DIODE(_02335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07283__A (.DIODE(_02259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07284__A (.DIODE(_02456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07284__B (.DIODE(_02467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07288__A1 (.DIODE(_00891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07288__A2 (.DIODE(_01000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07289__A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__07289__B (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__07289__C (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__07289__D (.DIODE(_00869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07290__A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__07290__B1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__07290__B2 (.DIODE(_00869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07292__A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__07292__B (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__07301__A (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__07302__A1 (.DIODE(_02664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07302__A2 (.DIODE(_00672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07303__B (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__07303__C (.DIODE(_00573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07303__D (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__07304__A2 (.DIODE(_00639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07304__B1 (.DIODE(_00573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07304__B2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__07306__A (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__07307__A (.DIODE(_01470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07307__B (.DIODE(_02719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07325__A1 (.DIODE(_00464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07325__A2 (.DIODE(_00530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07326__A (.DIODE(_00464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07326__B (.DIODE(_00530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07327__A1 (.DIODE(_00344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07327__A2 (.DIODE(_00410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07329__A (.DIODE(_02960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07330__A (.DIODE(_02971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07331__A (.DIODE(_02982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07332__A (.DIODE(_02993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07333__A (.DIODE(_03004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07334__A1 (.DIODE(_02138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07334__A2 (.DIODE(_00410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07334__B1 (.DIODE(_03015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07334__B2 (.DIODE(_00333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07335__A (.DIODE(_01470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07335__B (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__07335__C (.DIODE(_00355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07335__D (.DIODE(_02971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07337__A (.DIODE(_02018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07338__A (.DIODE(_03059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07339__A1 (.DIODE(_03070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07339__A2 (.DIODE(_02259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07339__B1 (.DIODE(_02171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07339__B2 (.DIODE(_02280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07340__A (.DIODE(_02007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07340__B (.DIODE(_02029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07340__C (.DIODE(_02105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07340__D (.DIODE(_02149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07344__A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__07344__A2 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__07345__A (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__07346__A1 (.DIODE(_01044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07346__A2 (.DIODE(_00880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07346__B1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__07347__A (.DIODE(_01044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07347__C (.DIODE(_00880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07347__D (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__07356__A (.DIODE(_02719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07357__A1 (.DIODE(_01744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07357__A2 (.DIODE(_03268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07358__A1 (.DIODE(_01295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07358__A2 (.DIODE(_02664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07358__B1 (.DIODE(_02719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07358__B2 (.DIODE(_01306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07359__A (.DIODE(_01295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07359__B (.DIODE(_01405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07359__C (.DIODE(_02664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07359__D (.DIODE(_02719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07372__A1 (.DIODE(_02456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07372__A2 (.DIODE(_02467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07377__A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__07378__A (.DIODE(_03499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07379__A (.DIODE(_03510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07380__A (.DIODE(_03521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07381__A (.DIODE(_03532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07382__A (.DIODE(_03543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07383__A1 (.DIODE(_00453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07383__A2 (.DIODE(_03554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07383__B1 (.DIODE(_00519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07383__B2 (.DIODE(_02051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07384__A (.DIODE(_00431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07385__A (.DIODE(_00978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07386__A (.DIODE(_03576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07386__B (.DIODE(_03587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07386__C (.DIODE(_03499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07386__D (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__07388__B (.DIODE(_03609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07394__A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__07395__A (.DIODE(_03685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07396__A (.DIODE(_03696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07397__A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__07398__A (.DIODE(_03718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07400__A (.DIODE(_02127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07400__B (.DIODE(_00322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07400__C (.DIODE(_03707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07400__D (.DIODE(_03740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07401__A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__07402__A (.DIODE(_03762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07403__A (.DIODE(_00322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07403__B (.DIODE(_03773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07404__B (.DIODE(_01470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07404__C (.DIODE(_03685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07404__D (.DIODE(_03718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07405__A2 (.DIODE(_03685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07405__B1 (.DIODE(_03718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07405__B2 (.DIODE(_01470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07409__A (.DIODE(_01197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07410__C (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__07410__D (.DIODE(_03718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07411__A2 (.DIODE(_03685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07411__B1 (.DIODE(_03718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07411__B2 (.DIODE(_01306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07413__A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__07414__A (.DIODE(_02127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07414__B (.DIODE(_03894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07416__A1 (.DIODE(_00311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07416__A2 (.DIODE(_03762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07417__A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__07418__A (.DIODE(_00311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07418__B (.DIODE(_03938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07424__A (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__07425__A (.DIODE(_04015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07426__A (.DIODE(_04026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07427__A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__07428__A (.DIODE(_04048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07429__A (.DIODE(_00442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07429__B (.DIODE(_02051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07429__C (.DIODE(_04037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07429__D (.DIODE(_04059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07430__A (.DIODE(_01284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07431__A (.DIODE(_04081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07431__B (.DIODE(_04048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07432__A (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__07433__A (.DIODE(_03576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07433__B (.DIODE(_03587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07433__C (.DIODE(_04015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07434__A1 (.DIODE(_03587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07434__A2 (.DIODE(_04015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07434__B2 (.DIODE(_03576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07438__A (.DIODE(_00978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07439__A (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__07440__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__07441__A (.DIODE(_00431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07441__B (.DIODE(_04169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07442__A1 (.DIODE(_03587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07442__B2 (.DIODE(_03576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07444__A (.DIODE(_01372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07444__B (.DIODE(_04026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07446__A1 (.DIODE(_01284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07446__A2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__07447__A (.DIODE(_01230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07448__A (.DIODE(_04268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07448__B (.DIODE(_04048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07454__A (.DIODE(_01996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07454__B (.DIODE(_00901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07454__C (.DIODE(_00366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07454__D (.DIODE(_02982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07455__A1 (.DIODE(_02018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07455__A2 (.DIODE(_00388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07455__B1 (.DIODE(_03004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07455__B2 (.DIODE(_02040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07457__A (.DIODE(_04367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07458__A1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__07458__A2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__07459__A (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__07459__C (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__07460__A1 (.DIODE(_01470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07460__A2 (.DIODE(_04378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07461__A (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__07462__A1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__07465__A (.DIODE(_00661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07467__A1 (.DIODE(_00661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07468__C (.DIODE(_04378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07469__A (.DIODE(_00573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07470__A1 (.DIODE(_01197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07470__A2 (.DIODE(_04367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07470__B2 (.DIODE(_04510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07478__A2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__07478__B2 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__07479__B (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__07479__C (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__07480__A1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__07480__A2 (.DIODE(_04367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07481__A (.DIODE(_00300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07481__B (.DIODE(_04598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07483__A (.DIODE(_00661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07483__B (.DIODE(_04367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07485__A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__07490__A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__07490__B (.DIODE(_04367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07500__A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__07501__A (.DIODE(_04851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07502__A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__07503__A (.DIODE(_01744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07503__B (.DIODE(_00311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07503__C (.DIODE(_04862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07503__D (.DIODE(_04873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07504__A (.DIODE(_04862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07505__A (.DIODE(_04895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07506__A (.DIODE(_04906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07507__A (.DIODE(_04873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07508__A (.DIODE(_04928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07509__A1 (.DIODE(_00333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07509__A2 (.DIODE(_04917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07509__B1 (.DIODE(_04939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07509__B2 (.DIODE(_02138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07513__A (.DIODE(_00573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07513__B (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__07513__C (.DIODE(_04851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07513__D (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__07514__A1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__07514__A2 (.DIODE(_04851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07514__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__07514__B2 (.DIODE(_00573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07516__A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__07517__A (.DIODE(_00300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07517__B (.DIODE(_05027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07522__B (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__07522__C (.DIODE(_00355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07522__D (.DIODE(_02960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07523__A2 (.DIODE(_00355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07523__B1 (.DIODE(_02960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07523__B2 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__07524__C (.DIODE(_00901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07524__D (.DIODE(_04378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07526__A1_N (.DIODE(_00901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07526__A2_N (.DIODE(_04378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07530__A (.DIODE(_04598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07531__A (.DIODE(_04378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07532__A (.DIODE(_05192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07533__A (.DIODE(_01405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07533__B (.DIODE(_05203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07534__A (.DIODE(_01361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07534__B (.DIODE(_05181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07541__B (.DIODE(_05291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07542__A (.DIODE(_00333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07542__B (.DIODE(_04939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07545__A (.DIODE(_02335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07545__B (.DIODE(_00399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07546__A1 (.DIODE(_02456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07546__A2 (.DIODE(_00399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07554__A (.DIODE(_01044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07555__A (.DIODE(_05445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07557__A (.DIODE(_05467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07558__A (.DIODE(_05478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07558__B (.DIODE(_01383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07559__A (.DIODE(_05456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07559__B (.DIODE(_01350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07565__A (.DIODE(_03268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07566__A (.DIODE(_02664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07567__A (.DIODE(_05577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07568__A (.DIODE(_01405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07568__B (.DIODE(_05588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07569__A (.DIODE(_01361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07569__B (.DIODE(_05566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07581__A (.DIODE(_00639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07582__A (.DIODE(_05731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07582__B (.DIODE(_01000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07582__C (.DIODE(_00628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07582__D (.DIODE(_05742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07583__A1 (.DIODE(_05731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07583__A2 (.DIODE(_00628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07583__B1 (.DIODE(_05742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07583__B2 (.DIODE(_01000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07584__C (.DIODE(_00901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07584__D (.DIODE(_02664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07586__A1_N (.DIODE(_02029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07586__A2_N (.DIODE(_05588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07589__A (.DIODE(_05445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07589__B (.DIODE(_05467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07589__C (.DIODE(_02105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07589__D (.DIODE(_00650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07590__A1 (.DIODE(_05456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07590__A2 (.DIODE(_02105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07590__B1 (.DIODE(_00650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07590__B2 (.DIODE(_05467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07592__A (.DIODE(_02007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07592__B (.DIODE(_05588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07594__B1 (.DIODE(_02029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07594__C1 (.DIODE(_05566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07595__A1 (.DIODE(_02029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07595__A2 (.DIODE(_05566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07623__A1 (.DIODE(_02007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07623__A2 (.DIODE(_05588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07624__A (.DIODE(_05445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07624__B (.DIODE(_05467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07624__C (.DIODE(_05742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07624__D (.DIODE(_02664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07625__A (.DIODE(_05467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07625__B (.DIODE(_00541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07626__A1 (.DIODE(_05445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07626__A2 (.DIODE(_00650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07627__C (.DIODE(_01996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07627__D (.DIODE(_03268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07628__A1_N (.DIODE(_02007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07628__A2_N (.DIODE(_05566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07644__A (.DIODE(_05456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07645__A (.DIODE(_06417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07646__A (.DIODE(_05478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07647__A (.DIODE(_06439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07648__A (.DIODE(_05588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07649__A (.DIODE(_06461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07650__A (.DIODE(_05566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07651__A (.DIODE(_06483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07652__A (.DIODE(_06428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07652__B (.DIODE(_06450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07652__C (.DIODE(_06472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07652__D (.DIODE(_06494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07653__A1 (.DIODE(_06428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07653__A2 (.DIODE(_06472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07653__B1 (.DIODE(_06483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07653__B2 (.DIODE(_06439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07663__A (.DIODE(_06428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07664__A (.DIODE(_06494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07665__A (.DIODE(_06626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07665__B (.DIODE(_06637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07673__A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__07674__A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__07675__A (.DIODE(_00442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07675__B (.DIODE(_00989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07675__C (.DIODE(_06733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07675__D (.DIODE(_06744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07676__A (.DIODE(_06733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07677__A (.DIODE(_06744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07678__A1 (.DIODE(_00442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07678__A2 (.DIODE(_06765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07678__B1 (.DIODE(_06775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07678__B2 (.DIODE(_02051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07680__A1 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07680__A2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__07680__B1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__07680__B2 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__07681__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07681__B (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__07681__C (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__07681__D (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__07682__A1 (.DIODE(_01076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07682__A2 (.DIODE(_03499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07683__A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__07683__B (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__07683__C (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__07683__D (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__07684__A1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__07684__A2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__07684__B1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__07684__B2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__07686__A (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__07686__B (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__07688__A1 (.DIODE(_01120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07688__A2 (.DIODE(_03499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07689__A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__07690__A (.DIODE(_06818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07691__A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__07692__A (.DIODE(_06820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07693__A (.DIODE(_00891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07693__B (.DIODE(_01120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07693__C (.DIODE(_06819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07693__D (.DIODE(_06821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07694__A1 (.DIODE(_01076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07694__A2 (.DIODE(_06818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07694__B1 (.DIODE(_06820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07694__B2 (.DIODE(_01120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07701__A1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__07701__A2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__07701__B1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__07701__B2 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07702__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07702__B (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__07702__C (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__07702__D (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__07703__A1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__07703__A2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__07704__A (.DIODE(_01230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07704__B (.DIODE(_00475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07706__A (.DIODE(_00880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07706__B (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__07708__A (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__07708__B (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__07713__A (.DIODE(_00880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07713__B (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__07723__A (.DIODE(_02105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07723__B (.DIODE(_00650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07723__C (.DIODE(_03510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07723__D (.DIODE(_00475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07724__A1 (.DIODE(_02259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07724__A2 (.DIODE(_03543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07724__B1 (.DIODE(_00508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07724__B2 (.DIODE(_02171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07728__A (.DIODE(_00563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07728__B (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__07728__C (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__07728__D (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__07729__A1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__07729__A2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__07729__B1 (.DIODE(_06820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07729__B2 (.DIODE(_00563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07731__A (.DIODE(_02664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07731__B (.DIODE(_00475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07736__A (.DIODE(_00420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07736__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__07736__C (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__07736__D (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__07737__A1 (.DIODE(_00420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07737__A2 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__07737__B1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__07737__B2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__07739__A (.DIODE(_01284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07739__B (.DIODE(_06744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07744__A (.DIODE(_06819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07745__A (.DIODE(_06821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07746__A (.DIODE(_06874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07747__A (.DIODE(_01383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07747__B (.DIODE(_06875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07748__A (.DIODE(_01350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07748__B (.DIODE(_06873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07755__A (.DIODE(_02259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07755__B (.DIODE(_00508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07756__A (.DIODE(_06775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07759__A (.DIODE(_00453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07759__B (.DIODE(_06885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07760__A1 (.DIODE(_00442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07760__A2 (.DIODE(_06775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07771__B (.DIODE(_00573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07771__C (.DIODE(_04851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07771__D (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__07772__A1 (.DIODE(_01208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07772__A2 (.DIODE(_04851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07772__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__07774__A (.DIODE(_01470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07774__B (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__07776__A1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__07776__A2 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__07777__A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__07777__B (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__07783__A (.DIODE(_01044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07783__C (.DIODE(_00355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07783__D (.DIODE(_02960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07784__A1 (.DIODE(_01044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07784__A2 (.DIODE(_00355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07784__B1 (.DIODE(_02960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07786__A (.DIODE(_01000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07786__B (.DIODE(_04378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07788__A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__07788__A2 (.DIODE(_04367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07789__A (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__07804__B (.DIODE(_05291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07808__A (.DIODE(_06472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07809__A (.DIODE(_06626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07809__B (.DIODE(_06450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07809__C (.DIODE(_06937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07809__D (.DIODE(_06637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07810__C1 (.DIODE(_06938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07811__A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__07811__B (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__07811__C (.DIODE(_06818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07811__D (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__07812__A1 (.DIODE(_00563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07812__A2 (.DIODE(_06818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07812__B1 (.DIODE(_06820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07812__B2 (.DIODE(_00639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07814__A (.DIODE(_00541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07814__B (.DIODE(_03499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07816__A1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__07816__A2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__07817__A (.DIODE(_02719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07817__B (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__07823__A (.DIODE(_00420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07823__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__07823__C (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__07823__D (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__07824__A1 (.DIODE(_00420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07824__A2 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__07824__B1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__07824__B2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__07826__A (.DIODE(_01076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07826__B (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__07828__A1 (.DIODE(_00880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07828__A2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__07829__A (.DIODE(_01120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07829__B (.DIODE(_06744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07835__A (.DIODE(_06873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07836__A (.DIODE(_06964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07837__A (.DIODE(_06875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07838__A (.DIODE(_01383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07838__B (.DIODE(_01350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07838__C (.DIODE(_06965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07838__D (.DIODE(_06966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07841__B (.DIODE(_06967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07842__A1 (.DIODE(_06967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07872__A (.DIODE(_00530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07872__B (.DIODE(_00410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07875__A (.DIODE(_06885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07876__A (.DIODE(_02467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07876__B (.DIODE(_07004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07878__A (.DIODE(_01230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07878__B (.DIODE(_06744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07880__A1 (.DIODE(_00891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07880__A2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__07881__A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__07882__A1 (.DIODE(_00978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07882__A2 (.DIODE(_07010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07882__B1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__07882__B2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__07883__A (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__07883__B (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__07883__C (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__07883__D (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__07885__A (.DIODE(_01120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07885__B (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__07890__A (.DIODE(_02719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07890__B (.DIODE(_00475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07892__A1 (.DIODE(_00541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07892__A2 (.DIODE(_03499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07893__A1 (.DIODE(_00639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07893__A2 (.DIODE(_06818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07893__B1 (.DIODE(_06820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07893__B2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__07894__A (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__07894__B (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__07894__C (.DIODE(_06818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07894__D (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__07896__A (.DIODE(_02719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07896__B (.DIODE(_03499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07911__A (.DIODE(_04939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07912__A (.DIODE(_02456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07912__B (.DIODE(_07040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07914__A (.DIODE(_00901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07916__A1 (.DIODE(_01996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07916__A2 (.DIODE(_04378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07917__A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__07917__B1 (.DIODE(_04367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07917__B2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__07918__A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__07918__B (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__07919__C (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__07920__A1_N (.DIODE(_01000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07929__A1 (.DIODE(_00672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07929__A2 (.DIODE(_05027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07930__A2 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__07930__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__07931__A (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__07931__C (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__07931__D (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__07932__C (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__07932__D (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__07933__A1_N (.DIODE(_01470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07933__A2_N (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__07947__B (.DIODE(_07075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07955__A (.DIODE(_03532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07955__B (.DIODE(_00497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07955__C (.DIODE(_00388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07955__D (.DIODE(_03004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07957__A1 (.DIODE(_03554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07957__A2 (.DIODE(_00410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07957__B1 (.DIODE(_03015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07957__B2 (.DIODE(_00519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07959__A (.DIODE(_06765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07960__A (.DIODE(_00003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07961__A1 (.DIODE(_02259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07961__A2 (.DIODE(_00004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07961__B1 (.DIODE(_07004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07961__B2 (.DIODE(_02171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07962__A (.DIODE(_02259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07962__B (.DIODE(_02171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07962__C (.DIODE(_00004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07962__D (.DIODE(_06885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07965__A1 (.DIODE(_01120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07965__A2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__07966__A1 (.DIODE(_01076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07966__A2 (.DIODE(_07010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07966__B1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__07966__B2 (.DIODE(_01120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07967__A (.DIODE(_00891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07967__B (.DIODE(_01120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07967__C (.DIODE(_07010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07967__D (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__07977__A1 (.DIODE(_02719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07977__A2 (.DIODE(_03499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07978__A1 (.DIODE(_00541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07978__A2 (.DIODE(_06818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07978__B1 (.DIODE(_06821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07978__B2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__07979__A (.DIODE(_00541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07979__B (.DIODE(_02719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07979__C (.DIODE(_06819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07979__D (.DIODE(_06821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07999__A1 (.DIODE(_02335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07999__A2 (.DIODE(_04917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07999__B1 (.DIODE(_04939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07999__B2 (.DIODE(_03070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08000__A (.DIODE(_03059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08000__B (.DIODE(_02040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08000__C (.DIODE(_04917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08000__D (.DIODE(_04939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08004__A1 (.DIODE(_01044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08004__A2 (.DIODE(_04367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08005__A (.DIODE(_01044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08005__C (.DIODE(_04367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08015__A1 (.DIODE(_01197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08015__A2 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__08015__B1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__08015__B2 (.DIODE(_01208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08016__A (.DIODE(_01197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08016__B (.DIODE(_04510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08016__C (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__08016__D (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__08034__B (.DIODE(_07075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08035__A2 (.DIODE(_07075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08042__A (.DIODE(_00002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08047__A (.DIODE(_03521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08047__B (.DIODE(_00377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08047__C (.DIODE(_02982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08047__D (.DIODE(_06875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08048__A1 (.DIODE(_03521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08048__A2 (.DIODE(_02993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08048__B1 (.DIODE(_06875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08048__B2 (.DIODE(_00377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08050__A (.DIODE(_05203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08051__A (.DIODE(_00094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08052__A (.DIODE(_00497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08052__B (.DIODE(_00095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08057__A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__08058__A (.DIODE(_00628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08058__B (.DIODE(_00650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08058__C (.DIODE(_00101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08058__D (.DIODE(_06733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08060__A1 (.DIODE(_02105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08060__A2 (.DIODE(_00101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08060__B1 (.DIODE(_06733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08060__B2 (.DIODE(_00650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08061__A (.DIODE(_05588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08061__B (.DIODE(_06744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08062__A1 (.DIODE(_06472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08062__A2 (.DIODE(_06885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08068__A (.DIODE(_07010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08069__A (.DIODE(_00112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08070__A (.DIODE(_00101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08071__A (.DIODE(_01383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08071__B (.DIODE(_00114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08072__A (.DIODE(_01350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08072__B (.DIODE(_00113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08077__A (.DIODE(_06874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08078__A (.DIODE(_06461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08078__B (.DIODE(_00121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08079__A (.DIODE(_05566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08079__B (.DIODE(_06964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08094__A (.DIODE(_05478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08095__A (.DIODE(_00138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08095__B (.DIODE(_02007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08095__C (.DIODE(_04928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08096__A1 (.DIODE(_02018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08096__A2 (.DIODE(_04895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08096__B1 (.DIODE(_04928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08096__B2 (.DIODE(_05478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08097__A1 (.DIODE(_04917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08098__A (.DIODE(_05027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08099__A (.DIODE(_00142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08100__A (.DIODE(_00143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08101__A (.DIODE(_00144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08102__A (.DIODE(_02280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08102__B (.DIODE(_00145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08107__A (.DIODE(_05181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08108__A (.DIODE(_05478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08108__B (.DIODE(_00094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08109__A (.DIODE(_06417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08109__B (.DIODE(_00151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08113__A (.DIODE(_01361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08114__A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__08115__A (.DIODE(_01405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08116__A (.DIODE(_00159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08116__B (.DIODE(_00142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08117__A (.DIODE(_00157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08117__B (.DIODE(_00158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08130__A2 (.DIODE(_07075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08132__B (.DIODE(_00175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08134__A (.DIODE(_00100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08135__B (.DIODE(_00002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08172__A (.DIODE(_00208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08178__A2 (.DIODE(_00219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08179__A2 (.DIODE(_00219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08181__A2 (.DIODE(_03609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08182__A2 (.DIODE(_03609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08183__B (.DIODE(_00219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08193__B1_N (.DIODE(_00208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08209__B1 (.DIODE(_00100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08210__B (.DIODE(_00175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08213__A (.DIODE(_00113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08214__A (.DIODE(_00114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08215__A (.DIODE(_01383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08215__B (.DIODE(_01350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08215__C (.DIODE(_00257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08215__D (.DIODE(_00258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08218__A (.DIODE(_06965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08219__A (.DIODE(_06966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08220__A (.DIODE(_06472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08220__B (.DIODE(_06483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08220__C (.DIODE(_00262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08220__D (.DIODE(_00263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08224__A (.DIODE(_00101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08225__A (.DIODE(_02116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08225__B (.DIODE(_02149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08225__C (.DIODE(_00112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08225__D (.DIODE(_00268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08226__A1 (.DIODE(_02116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08226__A2 (.DIODE(_00112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08226__B1 (.DIODE(_00268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08226__B2 (.DIODE(_02149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08228__A (.DIODE(_06461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08228__B (.DIODE(_00003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08231__A (.DIODE(_05566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08231__B (.DIODE(_06775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08249__A (.DIODE(_00095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08250__A (.DIODE(_00151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08251__A (.DIODE(_06428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08251__B (.DIODE(_06450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08251__C (.DIODE(_00293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08251__D (.DIODE(_00294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08254__A (.DIODE(_00158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08255__A (.DIODE(_00157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08255__B (.DIODE(_00159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08255__C (.DIODE(_00144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08255__D (.DIODE(_00298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08259__A (.DIODE(_06417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08259__B (.DIODE(_00138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08259__C (.DIODE(_04906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08259__D (.DIODE(_04928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08260__A1 (.DIODE(_00138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08260__A2 (.DIODE(_04906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08260__B1 (.DIODE(_04928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08260__B2 (.DIODE(_06417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08261__C (.DIODE(_02018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08261__D (.DIODE(_00143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08262__A1_N (.DIODE(_03059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08262__A2_N (.DIODE(_00144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08263__A1 (.DIODE(_02040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08263__A2 (.DIODE(_00143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08263__B2 (.DIODE(_04917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08264__A (.DIODE(_02040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08264__B (.DIODE(_00298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08265__A (.DIODE(_00298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08266__A1 (.DIODE(_02280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08266__A2 (.DIODE(_00310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08281__B (.DIODE(_00327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08283__A (.DIODE(_00377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08283__B (.DIODE(_02982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08283__C (.DIODE(_06873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08283__D (.DIODE(_06874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08284__A1 (.DIODE(_00377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08284__A2 (.DIODE(_06873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08284__B1 (.DIODE(_06875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08284__B2 (.DIODE(_02993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08286__A (.DIODE(_03532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08286__B (.DIODE(_00094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08288__A1 (.DIODE(_00497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08288__A2 (.DIODE(_00094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08289__A (.DIODE(_00497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08289__B (.DIODE(_00151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08295__B (.DIODE(_00342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08301__A (.DIODE(_04004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08318__A (.DIODE(_00354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08319__A (.DIODE(_00354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08320__A1 (.DIODE(_00352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08322__A (.DIODE(_04015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08323__A (.DIODE(_00373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08324__A (.DIODE(_00374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08326__A (.DIODE(_04059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08327__A (.DIODE(_00378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08328__A (.DIODE(_00379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08329__A (.DIODE(_00380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08330__A1 (.DIODE(_00464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08330__A2 (.DIODE(_00376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08330__B1 (.DIODE(_00381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08330__B2 (.DIODE(_02051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08332__A (.DIODE(_00383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08336__A (.DIODE(_03707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08337__A (.DIODE(_00389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08338__A (.DIODE(_00390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08339__A (.DIODE(_03740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08340__A (.DIODE(_00392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08341__A1 (.DIODE(_02138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08341__A2 (.DIODE(_00391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08341__B1 (.DIODE(_00393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08341__B2 (.DIODE(_00344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08343__B1 (.DIODE(_00395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08344__A (.DIODE(_00354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08345__A (.DIODE(_00352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08347__A (.DIODE(_00344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08347__B (.DIODE(_00391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08350__A (.DIODE(_00464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08350__B (.DIODE(_00381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08351__A1 (.DIODE(_00464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08351__A2 (.DIODE(_00381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08354__A (.DIODE(_00395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08359__A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__08360__A (.DIODE(_00413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08361__A (.DIODE(_00414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08362__A (.DIODE(_00415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08363__A (.DIODE(_00333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08363__B (.DIODE(_00416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08366__A1 (.DIODE(_02127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08366__A2 (.DIODE(_03894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08367__B (.DIODE(_04510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08367__C (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__08367__D (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__08368__A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__08369__A2 (.DIODE(_00423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08369__B1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__08369__B2 (.DIODE(_01306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08370__C (.DIODE(_00672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08370__D (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__08371__A1_N (.DIODE(_01744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08371__A2_N (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__08379__A (.DIODE(_02335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08379__B (.DIODE(_00389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08384__A (.DIODE(_02467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08384__B (.DIODE(_00381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08387__A1 (.DIODE(_04081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08387__A2 (.DIODE(_00373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08388__A (.DIODE(_00978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08388__B (.DIODE(_00880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08388__D (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__08389__A1 (.DIODE(_00880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08389__B2 (.DIODE(_04169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08391__A (.DIODE(_04268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08391__B (.DIODE(_04026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08399__A (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__08400__A (.DIODE(_00457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08401__A (.DIODE(_00458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08402__A (.DIODE(_00459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08403__A (.DIODE(_00453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08403__B (.DIODE(_00460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08407__B (.DIODE(_00327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08411__A1 (.DIODE(_06494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08411__A2 (.DIODE(_07004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08412__A1 (.DIODE(_02149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08412__A2 (.DIODE(_00112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08412__B1 (.DIODE(_00268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08412__B2 (.DIODE(_05588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08413__A (.DIODE(_02149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08413__B (.DIODE(_05577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08413__C (.DIODE(_07010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08413__D (.DIODE(_00101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08416__A (.DIODE(_06483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08416__B (.DIODE(_00003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08418__A1 (.DIODE(_06472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08418__A2 (.DIODE(_00003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08436__A (.DIODE(_05478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08436__B (.DIODE(_00142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08437__A1 (.DIODE(_05456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08437__A2 (.DIODE(_04895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08438__A (.DIODE(_05456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08438__B (.DIODE(_05478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08438__C (.DIODE(_00142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08438__D (.DIODE(_04862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08440__A (.DIODE(_02018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08440__B (.DIODE(_00158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08441__A1 (.DIODE(_03059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08441__A2 (.DIODE(_00158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08460__B (.DIODE(_00523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08462__A (.DIODE(_07040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08463__A (.DIODE(_00519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08463__B (.DIODE(_00526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08464__A (.DIODE(_00508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08464__B (.DIODE(_00294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08466__A1 (.DIODE(_03543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08466__A2 (.DIODE(_00095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08467__A (.DIODE(_02993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08467__B (.DIODE(_06873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08467__C (.DIODE(_06875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08467__D (.DIODE(_05203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08468__A1 (.DIODE(_02993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08468__A2 (.DIODE(_06873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08468__B1 (.DIODE(_06875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08468__B2 (.DIODE(_05203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08470__A (.DIODE(_03532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08470__B (.DIODE(_00151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08477__A (.DIODE(_07004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08478__A (.DIODE(_00543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08479__A (.DIODE(_00399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08479__B (.DIODE(_00544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08482__B (.DIODE(_00547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08483__B1_N (.DIODE(_00342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08495__A (.DIODE(_00439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08496__B1 (.DIODE(_04004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08504__A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__08505__A (.DIODE(_00571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08506__A (.DIODE(_00572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08507__A (.DIODE(_00574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08508__A1 (.DIODE(_02138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08508__A2 (.DIODE(_00415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08508__B1 (.DIODE(_00575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08508__B2 (.DIODE(_00333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08509__A (.DIODE(_01744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08509__B (.DIODE(_00311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08509__C (.DIODE(_00413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08509__D (.DIODE(_00571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08513__A1 (.DIODE(_01295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08513__A2 (.DIODE(_03894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08513__B1 (.DIODE(_03938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08513__B2 (.DIODE(_01405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08514__A (.DIODE(_01361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08514__B (.DIODE(_01405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08514__C (.DIODE(_03773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08514__D (.DIODE(_03938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08521__A1 (.DIODE(_03059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08521__A2 (.DIODE(_00389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08521__B1 (.DIODE(_00393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08521__B2 (.DIODE(_02280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08522__A (.DIODE(_02007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08522__B (.DIODE(_02040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08522__C (.DIODE(_03707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08522__D (.DIODE(_00392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08530__A1 (.DIODE(_00453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08530__A2 (.DIODE(_00460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08530__B1 (.DIODE(_02467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08530__B2 (.DIODE(_00380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08531__A1 (.DIODE(_02259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08531__A2 (.DIODE(_00376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08531__B1 (.DIODE(_00379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08531__B2 (.DIODE(_02171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08532__A (.DIODE(_02105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08532__B (.DIODE(_02149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08532__C (.DIODE(_04037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08532__D (.DIODE(_04048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08534__A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__08535__A (.DIODE(_00604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08536__A (.DIODE(_00605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08537__A (.DIODE(_00607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08538__A1 (.DIODE(_02051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08538__A2 (.DIODE(_00458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08538__B1 (.DIODE(_00608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08538__B2 (.DIODE(_00442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08539__A (.DIODE(_00453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08539__B (.DIODE(_02051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08539__C (.DIODE(_00458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08539__D (.DIODE(_00608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08540__A1 (.DIODE(_04268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08540__A2 (.DIODE(_04026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08543__A1 (.DIODE(_01230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08543__A2 (.DIODE(_00612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08543__B1 (.DIODE(_00613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08543__B2 (.DIODE(_01284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08544__A (.DIODE(_01372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08544__B (.DIODE(_04268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08544__C (.DIODE(_00612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08544__D (.DIODE(_00613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08559__A (.DIODE(_00410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08559__B (.DIODE(_00544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08562__A (.DIODE(_04917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08564__A1 (.DIODE(_00519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08564__A2 (.DIODE(_00636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08564__B1 (.DIODE(_00526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08564__B2 (.DIODE(_03554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08565__A (.DIODE(_03554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08565__B (.DIODE(_00508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08565__C (.DIODE(_04917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08565__D (.DIODE(_04939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08569__A1 (.DIODE(_03543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08569__A2 (.DIODE(_00294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08570__A1 (.DIODE(_06965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08570__A2 (.DIODE(_00293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08570__B1 (.DIODE(_00151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08570__B2 (.DIODE(_00263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08571__A (.DIODE(_06965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08571__B (.DIODE(_06966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08571__C (.DIODE(_00095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08571__D (.DIODE(_00151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08579__A (.DIODE(_00004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08580__A1 (.DIODE(_00399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08580__A2 (.DIODE(_00654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08580__B1 (.DIODE(_00543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08580__B2 (.DIODE(_03015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08581__A (.DIODE(_00388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08581__B (.DIODE(_02993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08581__C (.DIODE(_06765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08582__A (.DIODE(_00543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08591__B (.DIODE(_00523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08593__A1 (.DIODE(_06494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08593__A2 (.DIODE(_00004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08594__A (.DIODE(_00258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08595__A1 (.DIODE(_06472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08595__A2 (.DIODE(_00257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08595__B1 (.DIODE(_00670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08595__B2 (.DIODE(_06483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08596__A (.DIODE(_06472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08596__B (.DIODE(_06483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08596__C (.DIODE(_00113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08596__D (.DIODE(_00258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08611__A1 (.DIODE(_06428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08611__A2 (.DIODE(_00144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08611__B1 (.DIODE(_00310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08611__B2 (.DIODE(_06450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08612__A (.DIODE(_06428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08612__B (.DIODE(_06439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08612__C (.DIODE(_00144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08612__D (.DIODE(_00298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08625__B (.DIODE(_00703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08627__A (.DIODE(_00666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08628__B1 (.DIODE(_00547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08637__A (.DIODE(_00598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08638__A1 (.DIODE(_00439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08645__A (.DIODE(_00725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08649__A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__08650__A (.DIODE(_04510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08650__B (.DIODE(_00661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08650__C (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__08650__D (.DIODE(_00730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08651__A2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__08651__B1 (.DIODE(_00730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08651__B2 (.DIODE(_01470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08653__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__08654__A (.DIODE(_00311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08654__B (.DIODE(_00734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08659__A (.DIODE(_03938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08660__A (.DIODE(_03773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08661__A (.DIODE(_00159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08661__B (.DIODE(_00742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08662__A (.DIODE(_00157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08662__B (.DIODE(_00741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08663__A (.DIODE(_00741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08664__A1 (.DIODE(_00157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08664__A2 (.DIODE(_00745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08669__A (.DIODE(_05731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08669__B (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__08669__C (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__08669__D (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__08670__A1 (.DIODE(_05731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08670__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__08670__B1 (.DIODE(_03718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08670__B2 (.DIODE(_01000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08672__A (.DIODE(_03894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08673__A (.DIODE(_02029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08673__B (.DIODE(_00755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08683__A (.DIODE(_00563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08683__B (.DIODE(_00639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08683__C (.DIODE(_04015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08684__A1 (.DIODE(_00639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08684__A2 (.DIODE(_04015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08684__B2 (.DIODE(_00563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08686__A (.DIODE(_05577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08686__B (.DIODE(_04048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08692__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__08694__A (.DIODE(_00778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08697__A (.DIODE(_00782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08698__A (.DIODE(_00783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08699__A (.DIODE(_01383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08699__B (.DIODE(_00784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08700__A (.DIODE(_01350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08700__B (.DIODE(_00779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08704__A (.DIODE(_00442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08704__B (.DIODE(_00989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08704__C (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__08704__D (.DIODE(_00604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08705__A (.DIODE(_00431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08705__B (.DIODE(_04169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08705__C (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__08705__D (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__08706__A1 (.DIODE(_03587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08706__A2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__08706__B1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__08706__B2 (.DIODE(_00431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08708__A (.DIODE(_04081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08708__B (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__08719__A (.DIODE(_03532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08719__B (.DIODE(_00121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08719__C (.DIODE(_04895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08719__D (.DIODE(_04873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08720__A1 (.DIODE(_03532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08720__A2 (.DIODE(_04895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08720__B1 (.DIODE(_04873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08720__B2 (.DIODE(_00121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08721__C (.DIODE(_00497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08721__D (.DIODE(_00142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08723__A1_N (.DIODE(_00508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08723__A2_N (.DIODE(_00144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08729__A (.DIODE(_00294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08730__A (.DIODE(_00293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08731__A (.DIODE(_00263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08731__B (.DIODE(_00819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08732__A (.DIODE(_00262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08732__B (.DIODE(_00818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08736__A1 (.DIODE(_00377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08736__A2 (.DIODE(_00114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08736__B1 (.DIODE(_06765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08736__B2 (.DIODE(_02993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08737__A1 (.DIODE(_00258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08738__A (.DIODE(_06885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08738__B (.DIODE(_00293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08740__A (.DIODE(_07004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08741__A1 (.DIODE(_00543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08751__B (.DIODE(_00703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08752__A (.DIODE(_00257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08753__A (.DIODE(_00670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08754__A (.DIODE(_06937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08754__B (.DIODE(_00844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08755__A (.DIODE(_06637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08755__B (.DIODE(_00843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08756__C (.DIODE(_00846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08757__B1 (.DIODE(_00846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08766__A (.DIODE(_00310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08767__A (.DIODE(_06626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08767__B (.DIODE(_00859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08778__B (.DIODE(_00871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08781__B1_N (.DIODE(_00666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08794__A (.DIODE(_00765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08795__B1_N (.DIODE(_00598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08805__B (.DIODE(_04510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08805__C (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__08805__D (.DIODE(_00730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08806__A2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__08806__B1 (.DIODE(_00730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08808__A (.DIODE(_02127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08808__B (.DIODE(_00734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08810__A1 (.DIODE(_00300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08810__A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__08811__A (.DIODE(_00300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08811__B (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__08817__A (.DIODE(_00742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08818__A (.DIODE(_00914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08819__A (.DIODE(_00741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08820__A (.DIODE(_00157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08820__B (.DIODE(_00159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08820__C (.DIODE(_00915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08820__D (.DIODE(_00916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08822__A (.DIODE(_01044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08822__B (.DIODE(_05731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08822__C (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__08822__D (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__08823__A1 (.DIODE(_01044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08823__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__08823__B1 (.DIODE(_03718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08823__B2 (.DIODE(_05731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08825__A (.DIODE(_01996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08825__B (.DIODE(_03762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08827__A1 (.DIODE(_00901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08827__A2 (.DIODE(_03762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08828__A (.DIODE(_00901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08828__B (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__08845__A (.DIODE(_00563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08845__B (.DIODE(_00639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08846__A1 (.DIODE(_05742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08846__B2 (.DIODE(_00563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08848__A (.DIODE(_05577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08848__B (.DIODE(_04026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08850__A1 (.DIODE(_02664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08850__A2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__08851__A (.DIODE(_03268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08851__B (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__08857__A (.DIODE(_00431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08857__B (.DIODE(_04169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08857__C (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__08857__D (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__08858__A (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__08859__A1 (.DIODE(_03587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08859__A2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__08859__B1 (.DIODE(_00959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08859__B2 (.DIODE(_03576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08861__A (.DIODE(_01372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08861__B (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__08863__A1 (.DIODE(_01284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08863__A2 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__08864__A (.DIODE(_01230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08864__B (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__08889__A (.DIODE(_06965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08889__B (.DIODE(_06966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08889__C (.DIODE(_04906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08889__D (.DIODE(_04928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08890__A1 (.DIODE(_06966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08890__A2 (.DIODE(_04906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08890__B1 (.DIODE(_04928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08890__B2 (.DIODE(_06965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08892__A (.DIODE(_03543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08892__B (.DIODE(_00144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08894__B1 (.DIODE(_00508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08894__C1 (.DIODE(_00298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08895__A1 (.DIODE(_00508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08895__A2 (.DIODE(_00158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08903__A (.DIODE(_00377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08903__B (.DIODE(_02993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08903__C (.DIODE(_00112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08903__D (.DIODE(_00268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08904__A1 (.DIODE(_00388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08904__A2 (.DIODE(_00112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08904__B1 (.DIODE(_00114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08904__B2 (.DIODE(_03004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08905__C (.DIODE(_06765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08905__D (.DIODE(_00095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08906__A1_N (.DIODE(_00003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08906__A2_N (.DIODE(_00095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08908__A1 (.DIODE(_06775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08908__A2 (.DIODE(_00095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08908__B2 (.DIODE(_00258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08909__A (.DIODE(_06775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08909__B (.DIODE(_00151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08926__B (.DIODE(_00871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08932__B (.DIODE(_01039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08934__A (.DIODE(_01032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08939__A (.DIODE(_00991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08941__A (.DIODE(_00943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08942__A1 (.DIODE(_00765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08946__A (.DIODE(_00898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08948__A (.DIODE(_00410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08948__B (.DIODE(_00380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08949__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__08951__A (.DIODE(_01059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08952__A (.DIODE(_01060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08953__A (.DIODE(_01061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08956__A (.DIODE(_00460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08957__A (.DIODE(_02467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08957__B (.DIODE(_01066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08962__A1 (.DIODE(_04081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08962__A2 (.DIODE(_00604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08963__A (.DIODE(_04169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08963__B (.DIODE(_01076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08963__C (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__08963__D (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__08964__A1 (.DIODE(_01076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08964__A2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__08964__B1 (.DIODE(_00959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08964__B2 (.DIODE(_03587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08966__A (.DIODE(_04268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08966__B (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__08975__A1 (.DIODE(_05577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08975__A2 (.DIODE(_00373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08976__A (.DIODE(_00639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08976__B (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__08977__A1 (.DIODE(_00541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08977__B2 (.DIODE(_00639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08979__A (.DIODE(_03268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08979__B (.DIODE(_04026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08994__A (.DIODE(_00464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08994__B (.DIODE(_01062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08995__A (.DIODE(_01062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08996__A1 (.DIODE(_00464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08996__A2 (.DIODE(_01108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09000__B1_N (.DIODE(_01032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09001__B (.DIODE(_01039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09005__A (.DIODE(_06885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09005__B (.DIODE(_00294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09008__A1 (.DIODE(_03004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09008__A2 (.DIODE(_00113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09008__B1 (.DIODE(_00114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09008__B2 (.DIODE(_00095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09009__A (.DIODE(_03004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09009__B (.DIODE(_00113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09009__C (.DIODE(_00114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09009__D (.DIODE(_00094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09011__A (.DIODE(_00003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09011__B (.DIODE(_00151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09018__A1 (.DIODE(_03543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09018__A2 (.DIODE(_00144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09019__A (.DIODE(_06965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09019__B (.DIODE(_04906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09020__A (.DIODE(_06966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09020__B (.DIODE(_00142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09021__A (.DIODE(_06964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09021__B (.DIODE(_06966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09021__C (.DIODE(_00142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09021__D (.DIODE(_04895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09023__A1 (.DIODE(_03543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09023__A2 (.DIODE(_00298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09024__A (.DIODE(_03543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09024__B (.DIODE(_00298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09037__A (.DIODE(_00544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09038__A (.DIODE(_00526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09039__B1 (.DIODE(_01155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09039__C1 (.DIODE(_01156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09040__A1 (.DIODE(_01155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09040__A2 (.DIODE(_01156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09057__A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__09058__A (.DIODE(_01177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09059__A (.DIODE(_01178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09060__A (.DIODE(_01179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09061__A (.DIODE(_01180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09062__A (.DIODE(_01181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09063__A (.DIODE(_01182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09064__A (.DIODE(_00344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09064__B (.DIODE(_01183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09067__A (.DIODE(_00416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09068__A (.DIODE(_02456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09068__B (.DIODE(_01188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09072__A1 (.DIODE(_01996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09072__A2 (.DIODE(_03894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09073__A (.DIODE(_05445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09073__B (.DIODE(_05731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09073__C (.DIODE(_03718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09073__D (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__09074__A1 (.DIODE(_05445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09074__A2 (.DIODE(_00423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09074__B1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__09074__B2 (.DIODE(_05731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09075__C (.DIODE(_01996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09075__D (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__09076__A1_N (.DIODE(_01996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09076__A2_N (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__09085__A1 (.DIODE(_02127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09085__A2 (.DIODE(_00734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09086__C (.DIODE(_00730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09086__D (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__09087__A2 (.DIODE(_00730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09087__B1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__09087__B2 (.DIODE(_01306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09088__A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__09089__C (.DIODE(_01744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09089__D (.DIODE(_01211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09090__A1_N (.DIODE(_01744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09090__A2_N (.DIODE(_01211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09105__A (.DIODE(_00530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09105__B (.DIODE(_00391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09106__A1 (.DIODE(_00530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09106__A2 (.DIODE(_00391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09108__B (.DIODE(_01232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09109__B (.DIODE(_01233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09112__A1 (.DIODE(_00943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09119__A1 (.DIODE(_00344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09119__A2 (.DIODE(_01182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09121__A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__09124__A (.DIODE(_01248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09125__A (.DIODE(_01249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09126__A (.DIODE(_01250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09127__A1 (.DIODE(_02138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09127__A2 (.DIODE(_01182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09127__B1 (.DIODE(_01252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09127__B2 (.DIODE(_00344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09129__A (.DIODE(_02138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09129__B (.DIODE(_00322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09129__C (.DIODE(_01179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09129__D (.DIODE(_01254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09133__A1 (.DIODE(_05456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09133__A2 (.DIODE(_03773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09133__B1 (.DIODE(_03938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09133__B2 (.DIODE(_05467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09134__A (.DIODE(_03938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09135__A (.DIODE(_05456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09135__B (.DIODE(_05478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09135__C (.DIODE(_03773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09135__D (.DIODE(_01260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09145__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__09146__A1 (.DIODE(_01295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09146__A2 (.DIODE(_01272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09146__B1 (.DIODE(_01211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09146__B2 (.DIODE(_01405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09147__A (.DIODE(_01361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09147__B (.DIODE(_01405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09147__C (.DIODE(_01272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09147__D (.DIODE(_01211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09159__A (.DIODE(_00575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09160__A (.DIODE(_01288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09161__A1 (.DIODE(_03070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09161__A2 (.DIODE(_01188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09161__B1 (.DIODE(_01289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09161__B2 (.DIODE(_02456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09162__A (.DIODE(_03070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09162__B (.DIODE(_02280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09162__C (.DIODE(_00416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09162__D (.DIODE(_01288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09171__A1 (.DIODE(_03554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09171__A2 (.DIODE(_00391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09171__B1 (.DIODE(_00393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09171__B2 (.DIODE(_00519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09172__A (.DIODE(_03521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09172__B (.DIODE(_00486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09172__C (.DIODE(_03707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09172__D (.DIODE(_03740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09181__A (.DIODE(_00654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09182__A1 (.DIODE(_00544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09182__A2 (.DIODE(_00636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09182__B1 (.DIODE(_00526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09182__B2 (.DIODE(_01312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09183__A (.DIODE(_01312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09183__B (.DIODE(_00543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09183__C (.DIODE(_00636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09183__D (.DIODE(_00526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09188__A1 (.DIODE(_00257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09188__A2 (.DIODE(_00293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09188__B1 (.DIODE(_00294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09188__B2 (.DIODE(_00670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09189__A (.DIODE(_00257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09189__B (.DIODE(_00670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09189__C (.DIODE(_00819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09189__D (.DIODE(_00818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09200__A1 (.DIODE(_00262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09200__A2 (.DIODE(_00144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09200__B1 (.DIODE(_00298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09200__B2 (.DIODE(_00263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09201__A (.DIODE(_06965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09201__B (.DIODE(_06966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09201__C (.DIODE(_00143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09201__D (.DIODE(_00158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09210__B (.DIODE(_01343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09215__A1 (.DIODE(_01155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09215__A2 (.DIODE(_01156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09218__A (.DIODE(_01311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09218__B (.DIODE(_01352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09219__B_N (.DIODE(_01352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09223__A1 (.DIODE(_00991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09226__A1 (.DIODE(_00410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09226__A2 (.DIODE(_00376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09226__B1 (.DIODE(_00380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09226__B2 (.DIODE(_03015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09227__A (.DIODE(_00355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09227__B (.DIODE(_02960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09227__C (.DIODE(_04015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09228__A (.DIODE(_04048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09231__A1 (.DIODE(_01339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09231__A2 (.DIODE(_00604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09232__A (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__09233__A (.DIODE(_00959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09234__A1 (.DIODE(_04268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09234__A2 (.DIODE(_01368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09234__B1 (.DIODE(_01369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09234__B2 (.DIODE(_01372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09235__A (.DIODE(_01284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09235__B (.DIODE(_01230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09235__C (.DIODE(_01368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09235__D (.DIODE(_00959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09245__A1 (.DIODE(_05566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09245__A2 (.DIODE(_00373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09246__A1 (.DIODE(_03268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09246__A2 (.DIODE(_00612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09246__B1 (.DIODE(_00613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09246__B2 (.DIODE(_05577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09247__A (.DIODE(_02664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09247__B (.DIODE(_02719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09260__A (.DIODE(_02116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09260__C (.DIODE(_00605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09261__A (.DIODE(_00608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09262__A1 (.DIODE(_02171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09262__A2 (.DIODE(_00460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09262__B1 (.DIODE(_01400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09262__B2 (.DIODE(_02467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09263__A1 (.DIODE(_01066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09270__A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__09271__A (.DIODE(_01410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09272__A (.DIODE(_01411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09273__A (.DIODE(_01412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09274__A (.DIODE(_01413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09275__A (.DIODE(_01414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09276__A1 (.DIODE(_02051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09276__A2 (.DIODE(_01062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09276__B1 (.DIODE(_01415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09276__B2 (.DIODE(_00464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09277__A (.DIODE(_00431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09277__B (.DIODE(_04169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09277__C (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__09286__A (.DIODE(_01309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09289__A2 (.DIODE(_01233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09295__A1 (.DIODE(_00898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09304__A_N (.DIODE(_01311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09304__B (.DIODE(_01352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09305__B (.DIODE(_01343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09308__A (.DIODE(_00844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09308__B (.DIODE(_00819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09309__A (.DIODE(_00843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09309__B (.DIODE(_00818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09315__A (.DIODE(_00262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09315__B (.DIODE(_00859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09320__B (.DIODE(_01463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09324__A (.DIODE(_00844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09324__B (.DIODE(_00654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09325__A1 (.DIODE(_00654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09325__B1 (.DIODE(_07040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09325__B2 (.DIODE(_00844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09326__A1 (.DIODE(_00526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09327__A (.DIODE(_00145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09328__A (.DIODE(_01472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09329__A (.DIODE(_00544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09329__B (.DIODE(_01473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09341__B1 (.DIODE(_01486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09344__C_N (.DIODE(_01486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09347__A1 (.DIODE(_02960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09347__A2 (.DIODE(_04015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09347__B2 (.DIODE(_00355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09348__A1 (.DIODE(_00612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09349__A (.DIODE(_05192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09349__B (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__09356__A (.DIODE(_01369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09357__A (.DIODE(_01504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09358__A (.DIODE(_01368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09360__A (.DIODE(_01507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09361__A (.DIODE(_01383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09361__B (.DIODE(_01508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09362__A (.DIODE(_01350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09362__B (.DIODE(_01505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09368__A (.DIODE(_00779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09369__A (.DIODE(_00784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09370__A (.DIODE(_06461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09370__B (.DIODE(_01518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09371__A (.DIODE(_06483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09371__B (.DIODE(_01517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09380__A2 (.DIODE(_00605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09380__B1 (.DIODE(_01508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09380__B2 (.DIODE(_02116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09381__A (.DIODE(_01508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09383__A (.DIODE(_06472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09383__B (.DIODE(_00458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09385__A (.DIODE(_00459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09386__A1 (.DIODE(_00460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09394__A (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__09396__A1 (.DIODE(_04169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09396__A2 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__09396__B2 (.DIODE(_00431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09398__A (.DIODE(_01372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09398__B (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__09404__A (.DIODE(_01500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09411__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__09412__A1 (.DIODE(_04510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09412__A2 (.DIODE(_01177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09412__B2 (.DIODE(_00661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09414__A (.DIODE(_04510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09414__B (.DIODE(_00661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09414__C (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__09414__D (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__09415__A1_N (.DIODE(_00322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09415__A2_N (.DIODE(_01564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09416__B (.DIODE(_01564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09416__C (.DIODE(_00311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09421__A (.DIODE(_00138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09421__B (.DIODE(_00742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09422__A (.DIODE(_06428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09422__B (.DIODE(_00745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09423__A1 (.DIODE(_06417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09423__A2 (.DIODE(_00745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09429__A (.DIODE(_01211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09430__A (.DIODE(_01584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09431__A (.DIODE(_01272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09432__A (.DIODE(_00159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09432__B (.DIODE(_01586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09433__A (.DIODE(_00157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09433__B (.DIODE(_01585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09434__A1 (.DIODE(_00157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09434__A2 (.DIODE(_01584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09441__A (.DIODE(_06439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09441__B (.DIODE(_02018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09441__C (.DIODE(_00574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09442__A1 (.DIODE(_06439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09442__A2 (.DIODE(_00414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09442__B1 (.DIODE(_00574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09442__B2 (.DIODE(_02018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09443__A1 (.DIODE(_00416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09444__A (.DIODE(_01586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09445__A (.DIODE(_01600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09446__A (.DIODE(_02335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09446__B (.DIODE(_01601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09457__A1 (.DIODE(_06820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09457__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__09457__B1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__09457__B2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__09459__A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__09459__B (.DIODE(_06820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09459__C (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__09459__D (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__09460__A1_N (.DIODE(_00475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09460__A2_N (.DIODE(_03894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09461__B (.DIODE(_03894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09461__C (.DIODE(_00475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09468__B1 (.DIODE(_01626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09469__A (.DIODE(_01626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09471__B1 (.DIODE(_01309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09488__B (.DIODE(_00898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09490__A1 (.DIODE(_03587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09490__B1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__09490__B2 (.DIODE(_03576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09491__A (.DIODE(_00431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09491__B (.DIODE(_04169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09491__C (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__09491__D (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__09493__A (.DIODE(_01372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09493__B (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__09495__A (.DIODE(_00431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09495__B (.DIODE(_04169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09495__C (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__09495__D (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__09496__A1 (.DIODE(_01284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09496__A2 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__09497__A (.DIODE(_04268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09497__B (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__09503__A (.DIODE(_01508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09504__A2 (.DIODE(_01664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09504__B1 (.DIODE(_01505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09504__B2 (.DIODE(_02116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09505__A (.DIODE(_02116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09505__C (.DIODE(_01508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09505__D (.DIODE(_01504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09507__A (.DIODE(_06472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09507__B (.DIODE(_00607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09510__A (.DIODE(_06494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09510__B (.DIODE(_00458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09511__A1 (.DIODE(_06494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09511__A2 (.DIODE(_00459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09534__A1 (.DIODE(_02971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09534__B2 (.DIODE(_00366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09535__A (.DIODE(_00355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09535__B (.DIODE(_02960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09537__A (.DIODE(_05192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09537__B (.DIODE(_04026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09539__A (.DIODE(_00355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09539__B (.DIODE(_02960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09539__C (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__09540__A1 (.DIODE(_05192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09540__A2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__09541__A (.DIODE(_04598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09541__B (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__09547__B (.DIODE(_01712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09548__B1 (.DIODE(_01500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09557__A (.DIODE(_00843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09557__B (.DIODE(_00844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09557__D (.DIODE(_07040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09558__A1 (.DIODE(_00844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09558__B1 (.DIODE(_07040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09558__B2 (.DIODE(_00843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09559__C (.DIODE(_00654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09559__D (.DIODE(_01472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09560__A1_N (.DIODE(_00654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09560__A2_N (.DIODE(_01472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09561__A1 (.DIODE(_00543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09561__A2 (.DIODE(_01472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09561__B2 (.DIODE(_07040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09562__A (.DIODE(_00543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09562__B (.DIODE(_00859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09563__A1 (.DIODE(_00544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09563__A2 (.DIODE(_00859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09570__B (.DIODE(_01463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09574__B (.DIODE(_01741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09584__A (.DIODE(_01486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09584__B_N (.DIODE(_01752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09586__B (.DIODE(_01486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09587__A2_N (.DIODE(_01486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09588__A1 (.DIODE(_00991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09588__C1 (.DIODE(_01752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09591__A (.DIODE(_06818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09591__B (.DIODE(_06820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09591__C (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__09592__A1 (.DIODE(_06818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09592__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__09592__B1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__09592__B2 (.DIODE(_06820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09593__A1 (.DIODE(_03685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09594__A (.DIODE(_03510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09594__B (.DIODE(_03762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09596__A1 (.DIODE(_00475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09596__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__09597__A (.DIODE(_00475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09597__B (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__09603__A1 (.DIODE(_06428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09603__A2 (.DIODE(_00415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09603__B1 (.DIODE(_00574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09603__B2 (.DIODE(_06439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09604__A (.DIODE(_06417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09604__B (.DIODE(_00138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09604__C (.DIODE(_00414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09604__D (.DIODE(_00574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09606__A (.DIODE(_03059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09606__B (.DIODE(_01600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09608__A (.DIODE(_01585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09609__A1 (.DIODE(_02040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09609__A2 (.DIODE(_01600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09609__B2 (.DIODE(_00415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09610__A (.DIODE(_02280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09610__B (.DIODE(_01780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09611__A1 (.DIODE(_02335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09611__A2 (.DIODE(_01780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09634__A (.DIODE(_01197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09634__B (.DIODE(_04510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09634__C (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__09635__A1 (.DIODE(_01197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09635__A2 (.DIODE(_01177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09635__B2 (.DIODE(_04510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09636__A1 (.DIODE(_01177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09637__A (.DIODE(_01744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09637__B (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__09639__A1 (.DIODE(_00300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09639__A2 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__09640__A (.DIODE(_00311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09640__B (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__09653__C_N (.DIODE(_01828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09654__B1_N (.DIODE(_01828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09655__A1 (.DIODE(_01626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09662__B (.DIODE(_01741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09663__A (.DIODE(_00670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09663__B (.DIODE(_00145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09664__A1 (.DIODE(_00843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09665__A (.DIODE(_00843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09665__B (.DIODE(_00670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09665__C (.DIODE(_00145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09665__D (.DIODE(_04917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09667__A (.DIODE(_00654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09667__B (.DIODE(_00859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09668__A1 (.DIODE(_00654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09668__A2 (.DIODE(_00859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09689__B (.DIODE(_01867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09690__A (.DIODE(_04939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09690__B (.DIODE(_00379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09691__A (.DIODE(_05181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09691__B (.DIODE(_04059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09693__A1 (.DIODE(_05192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09693__A2 (.DIODE(_00373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09694__A1 (.DIODE(_04378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09694__B2 (.DIODE(_02971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09695__A (.DIODE(_02960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09695__B (.DIODE(_04367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09697__A (.DIODE(_04598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09697__B (.DIODE(_04026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09704__A (.DIODE(_00388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09704__B (.DIODE(_00459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09711__A1 (.DIODE(_06461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09711__A2 (.DIODE(_01508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09711__B1 (.DIODE(_01505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09712__B (.DIODE(_06461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09712__C (.DIODE(_01508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09712__D (.DIODE(_01504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09714__A1 (.DIODE(_06494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09714__A2 (.DIODE(_00608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09715__A (.DIODE(_06483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09715__B (.DIODE(_00607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09734__A (.DIODE(_02467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09734__B (.DIODE(_01060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09735__A (.DIODE(_01339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09737__A1 (.DIODE(_04081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09737__A2 (.DIODE(_01410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09738__A1 (.DIODE(_00891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09738__B1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__09738__B2 (.DIODE(_03587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09739__A (.DIODE(_04169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09739__B (.DIODE(_01076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09739__D (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__09741__A (.DIODE(_04268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09741__B (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__09748__A (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__09749__A (.DIODE(_01933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09750__A (.DIODE(_00453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09750__B (.DIODE(_01934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09756__A (.DIODE(_01889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09757__B1 (.DIODE(_01712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09766__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__09767__A (.DIODE(_01953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09768__A (.DIODE(_01954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09769__A (.DIODE(_01955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09770__A (.DIODE(_01956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09771__A (.DIODE(_01957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09772__A (.DIODE(_00344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09772__B (.DIODE(_01958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09773__A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__09774__A (.DIODE(_00322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09774__B (.DIODE(_01960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09776__A1_N (.DIODE(_01178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09777__A (.DIODE(_01295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09778__A (.DIODE(_01306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09778__B (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__09779__A (.DIODE(_01197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09779__B (.DIODE(_04510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09779__D (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__09781__A (.DIODE(_01744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09781__B (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__09788__A (.DIODE(_02456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09788__B (.DIODE(_01180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09789__A1 (.DIODE(_02456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09789__A2 (.DIODE(_01181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09794__A1 (.DIODE(_06417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09794__A2 (.DIODE(_00574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09794__B1 (.DIODE(_01600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09794__B2 (.DIODE(_06439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09795__A (.DIODE(_05456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09795__B (.DIODE(_00138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09795__C (.DIODE(_00572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09795__D (.DIODE(_01586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09797__A1 (.DIODE(_03070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09797__A2 (.DIODE(_01585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09798__A (.DIODE(_03059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09798__B (.DIODE(_01585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09816__A (.DIODE(_01188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09817__A (.DIODE(_00530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09817__B (.DIODE(_02008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09818__A (.DIODE(_00486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09818__B (.DIODE(_01260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09820__A1_N (.DIODE(_03696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09821__A (.DIODE(_06819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09821__B (.DIODE(_00423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09822__A (.DIODE(_06821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09822__B (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__09823__A (.DIODE(_06818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09823__B (.DIODE(_06820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09823__C (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__09823__D (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__09825__A (.DIODE(_03510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09825__B (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__09832__A (.DIODE(_07004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09832__B (.DIODE(_00390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09833__A1 (.DIODE(_07004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09833__A2 (.DIODE(_00390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09846__B (.DIODE(_02039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09847__A (.DIODE(_01828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09860__A2 (.DIODE(_02039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09862__A1 (.DIODE(_00519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09862__A2 (.DIODE(_01188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09864__A1 (.DIODE(_00004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09864__A2 (.DIODE(_00390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09864__B1 (.DIODE(_00393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09864__B2 (.DIODE(_07004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09865__A (.DIODE(_06765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09865__B (.DIODE(_06775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09865__C (.DIODE(_03707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09865__D (.DIODE(_03740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09867__A1 (.DIODE(_03521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09867__A2 (.DIODE(_01260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09868__A1 (.DIODE(_06873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09868__A2 (.DIODE(_00755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09868__B1 (.DIODE(_01260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09868__B2 (.DIODE(_06875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09869__A (.DIODE(_06964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09869__B (.DIODE(_00121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09869__C (.DIODE(_00755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09869__D (.DIODE(_00741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09880__A1 (.DIODE(_03554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09880__A2 (.DIODE(_00416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09880__B1 (.DIODE(_01288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09880__B2 (.DIODE(_00508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09881__A (.DIODE(_03521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09881__B (.DIODE(_00486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09881__C (.DIODE(_00413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09881__D (.DIODE(_00572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09890__A (.DIODE(_01780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09891__A1 (.DIODE(_03070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09891__A2 (.DIODE(_02088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09892__A (.DIODE(_01601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09893__A1 (.DIODE(_06626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09893__A2 (.DIODE(_02090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09893__B1 (.DIODE(_02088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09893__B2 (.DIODE(_06450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09894__A (.DIODE(_06626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09894__B (.DIODE(_06450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09894__C (.DIODE(_02090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09894__D (.DIODE(_02088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09910__A1 (.DIODE(_00333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09910__A2 (.DIODE(_01955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09912__A1 (.DIODE(_03070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09912__A2 (.DIODE(_01180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09912__B1 (.DIODE(_01249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09912__B2 (.DIODE(_02335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09913__A (.DIODE(_02007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09913__B (.DIODE(_02040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09913__C (.DIODE(_01179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09913__D (.DIODE(_01254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09915__A1 (.DIODE(_02138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09915__A2 (.DIODE(_01960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09916__A (.DIODE(_01564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09917__A1 (.DIODE(_01361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09917__A2 (.DIODE(_02117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09917__B1 (.DIODE(_01960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09917__B2 (.DIODE(_00159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09918__A (.DIODE(_02117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09919__A (.DIODE(_01960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09920__A (.DIODE(_01361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09920__B (.DIODE(_00159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09920__C (.DIODE(_02119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09920__D (.DIODE(_02120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09931__A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__09932__A (.DIODE(_02133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09933__A (.DIODE(_02134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09934__A1 (.DIODE(_02138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09934__A2 (.DIODE(_01954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09934__B1 (.DIODE(_02135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09934__B2 (.DIODE(_00333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09935__A (.DIODE(_02127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09935__B (.DIODE(_00322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09935__C (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__09935__D (.DIODE(_02133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09947__B1 (.DIODE(_02150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09951__A1 (.DIODE(_01339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09951__A2 (.DIODE(_01410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09952__A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__09953__A1 (.DIODE(_04268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09953__B2 (.DIODE(_01372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09955__A (.DIODE(_04081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09955__B (.DIODE(_01339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09955__C (.DIODE(_02158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09963__A (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__09964__A (.DIODE(_02168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09965__A1 (.DIODE(_02051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09965__A2 (.DIODE(_01934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09965__B1 (.DIODE(_02169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09965__B2 (.DIODE(_00453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09966__A (.DIODE(_03576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09966__B (.DIODE(_00989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09966__C (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__09967__A (.DIODE(_01934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09970__A1 (.DIODE(_02171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09970__A2 (.DIODE(_01060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09970__B1 (.DIODE(_01413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09970__B2 (.DIODE(_02259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09971__A (.DIODE(_02105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09971__B (.DIODE(_02149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09971__D (.DIODE(_01411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09979__A1 (.DIODE(_06637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09979__A2 (.DIODE(_01400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09980__A (.DIODE(_01664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09981__A (.DIODE(_02187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09982__A (.DIODE(_01505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09983__A (.DIODE(_02189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09984__A1 (.DIODE(_06637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09984__A2 (.DIODE(_02188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09984__B1 (.DIODE(_02190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09984__B2 (.DIODE(_06937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09985__A (.DIODE(_06937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09985__B (.DIODE(_06637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09985__C (.DIODE(_02187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09985__D (.DIODE(_02189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10003__A1 (.DIODE(_05181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10003__A2 (.DIODE(_04037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10004__A1 (.DIODE(_04598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10004__A2 (.DIODE(_00612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10004__B1 (.DIODE(_00613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10004__B2 (.DIODE(_05192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10005__A (.DIODE(_05203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10005__B (.DIODE(_04598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10005__C (.DIODE(_00782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10005__D (.DIODE(_00613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10013__A1 (.DIODE(_03015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10013__A2 (.DIODE(_00458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10013__B1 (.DIODE(_00608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10013__B2 (.DIODE(_00388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10014__A (.DIODE(_00366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10014__B (.DIODE(_02971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10014__C (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__10015__A (.DIODE(_00459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10018__A1 (.DIODE(_04939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10018__A2 (.DIODE(_00376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10018__B1 (.DIODE(_00379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10018__B2 (.DIODE(_04917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10019__A (.DIODE(_04862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10019__B (.DIODE(_04873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10019__C (.DIODE(_04037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10019__D (.DIODE(_04059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10025__B (.DIODE(_02235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10026__B1 (.DIODE(_01889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10032__C1 (.DIODE(_01867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10034__A (.DIODE(_00843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10035__A (.DIODE(_00859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10036__A (.DIODE(_00844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10037__A1 (.DIODE(_02246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10037__A2 (.DIODE(_01473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10037__B1 (.DIODE(_02247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10037__B2 (.DIODE(_02249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10038__A (.DIODE(_02246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10038__B (.DIODE(_02249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10038__C (.DIODE(_01473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10038__D (.DIODE(_02247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10057__A (.DIODE(_02151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10064__B (.DIODE(_02278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10066__A (.DIODE(_01752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10066__B (.DIODE(_01867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10068__A (.DIODE(_02246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10068__B (.DIODE(_02247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10078__B (.DIODE(_02293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10079__B (.DIODE(_02293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10080__D1 (.DIODE(_01486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10081__A (.DIODE(_02293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10082__A1 (.DIODE(_00991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10088__A (.DIODE(_02304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10089__A (.DIODE(_02158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10090__A (.DIODE(_01383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10090__B (.DIODE(_02306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10091__A (.DIODE(_01350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10091__B (.DIODE(_02305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10092__B (.DIODE(_02308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10095__A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__10096__A1 (.DIODE(_00989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10096__A2 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__10096__B2 (.DIODE(_03576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10098__A (.DIODE(_04081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10098__B (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__10100__A (.DIODE(_01933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10101__A1 (.DIODE(_01934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10104__A1 (.DIODE(_00650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10104__A2 (.DIODE(_01410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10104__B1 (.DIODE(_02158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10104__B2 (.DIODE(_02105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10105__A (.DIODE(_00628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10105__B (.DIODE(_05742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10105__C (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__10106__A1_N (.DIODE(_05588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10107__A1 (.DIODE(_05742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10107__A2 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__10107__B2 (.DIODE(_00628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10108__C (.DIODE(_05577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10117__A (.DIODE(_06937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10117__B (.DIODE(_02188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10118__A (.DIODE(_06637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10118__B (.DIODE(_02190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10130__A (.DIODE(_00094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10130__B (.DIODE(_00784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10131__A (.DIODE(_00151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10131__B (.DIODE(_01517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10135__A1 (.DIODE(_02971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10135__A2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__10135__B1 (.DIODE(_01368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10135__B2 (.DIODE(_00366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10137__A (.DIODE(_05203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10137__B (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__10139__A (.DIODE(_00457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10140__A1 (.DIODE(_00458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10143__A1 (.DIODE(_04862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10143__A2 (.DIODE(_00373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10143__B1 (.DIODE(_00782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10143__B2 (.DIODE(_04873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10144__A (.DIODE(_04851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10144__B (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__10144__C (.DIODE(_04015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10145__A1_N (.DIODE(_05027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10145__A2_N (.DIODE(_04048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10146__A1 (.DIODE(_04851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10146__A2 (.DIODE(_04015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10146__B2 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__10147__B (.DIODE(_04048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10147__C (.DIODE(_05027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10155__B (.DIODE(_02377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10156__B1_N (.DIODE(_02235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10169__A (.DIODE(_06965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10169__B (.DIODE(_00741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10175__A1 (.DIODE(_00101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10175__A2 (.DIODE(_03685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10175__B1 (.DIODE(_03718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10175__B2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__10177__A (.DIODE(_00101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10177__B (.DIODE(_06733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10177__C (.DIODE(_03685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10177__D (.DIODE(_00423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10178__A1_N (.DIODE(_06744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10178__A2_N (.DIODE(_03773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10179__B (.DIODE(_03894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10179__C (.DIODE(_06744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10185__A1 (.DIODE(_06821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10185__A2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__10185__B1 (.DIODE(_00730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10185__B2 (.DIODE(_03499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10187__A (.DIODE(_03499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10187__B (.DIODE(_06821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10187__C (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__10187__D (.DIODE(_00730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10188__A1_N (.DIODE(_00486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10188__A2_N (.DIODE(_00734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10189__B (.DIODE(_00734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10189__C (.DIODE(_00486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10198__A (.DIODE(_02088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10199__A (.DIODE(_02090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10200__A (.DIODE(_06450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10200__B (.DIODE(_02427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10201__A (.DIODE(_06626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10201__B (.DIODE(_02426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10212__A (.DIODE(_00157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10212__B (.DIODE(_02120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10218__A1 (.DIODE(_05731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10218__A2 (.DIODE(_01177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10218__B2 (.DIODE(_01000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10220__A (.DIODE(_05467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10220__B (.DIODE(_01000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10220__C (.DIODE(_01177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10221__A1_N (.DIODE(_02029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10221__A2_N (.DIODE(_01564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10222__B (.DIODE(_01564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10222__C (.DIODE(_02029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10228__A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__10229__A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__10229__B1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__10229__B2 (.DIODE(_01470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10231__A (.DIODE(_01306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10231__B (.DIODE(_00672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10231__C (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__10231__D (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__10232__A1_N (.DIODE(_00322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10232__A2_N (.DIODE(_02459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10233__B (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__10233__C (.DIODE(_00322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10247__A2 (.DIODE(_02150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10248__B (.DIODE(_02150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10250__B1 (.DIODE(_02482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10251__C (.DIODE(_02482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10253__B1 (.DIODE(_02151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10265__A1 (.DIODE(_00991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10271__B (.DIODE(_02308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10273__A (.DIODE(_03576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10273__B (.DIODE(_00989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10274__A1 (.DIODE(_00989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10274__B1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__10274__B2 (.DIODE(_03576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10275__A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__10276__A (.DIODE(_04081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10276__B (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__10278__A1 (.DIODE(_01372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10278__A2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__10279__A (.DIODE(_01339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10279__B (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__10288__A (.DIODE(_00628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10288__B (.DIODE(_05742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10289__A1 (.DIODE(_05742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10289__B2 (.DIODE(_00628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10291__A (.DIODE(_05577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10291__B (.DIODE(_01410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10293__A1 (.DIODE(_05577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10293__A2 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__10294__A (.DIODE(_03268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10310__A (.DIODE(_00366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10310__B (.DIODE(_02971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10310__C (.DIODE(_01368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10311__A1 (.DIODE(_02971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10311__A2 (.DIODE(_01368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10311__B1 (.DIODE(_00959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10311__B2 (.DIODE(_00366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10312__A1 (.DIODE(_01369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10313__A (.DIODE(_05203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10313__B (.DIODE(_00604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10315__A1 (.DIODE(_05192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10315__A2 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__10316__A (.DIODE(_04598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10316__B (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__10325__A (.DIODE(_04862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10325__B (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__10326__A1 (.DIODE(_04851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10326__B2 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__10327__A1 (.DIODE(_00613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10328__A (.DIODE(_05027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10328__B (.DIODE(_00373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10330__A1 (.DIODE(_05027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10330__A2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__10331__A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__10331__B (.DIODE(_04048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10342__B (.DIODE(_02582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10345__A2 (.DIODE(_02377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10350__A1 (.DIODE(_02496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10350__A2 (.DIODE(_02498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10351__A (.DIODE(_02496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10351__B (.DIODE(_02498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10357__A (.DIODE(_07010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10357__B (.DIODE(_00101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10357__C (.DIODE(_00423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10358__A1 (.DIODE(_07010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10358__A2 (.DIODE(_03685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10358__B1 (.DIODE(_00423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10358__B2 (.DIODE(_00101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10359__A1 (.DIODE(_03696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10360__A (.DIODE(_06733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10360__B (.DIODE(_03773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10362__A1 (.DIODE(_06744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10362__A2 (.DIODE(_03894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10363__A (.DIODE(_06744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10363__B (.DIODE(_03938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10374__A (.DIODE(_06819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10374__B (.DIODE(_06821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10374__C (.DIODE(_00730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10375__A1 (.DIODE(_06819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10375__A2 (.DIODE(_00413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10375__B1 (.DIODE(_00571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10375__B2 (.DIODE(_06821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10376__A1 (.DIODE(_00413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10377__A (.DIODE(_03521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10377__B (.DIODE(_00734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10379__A1 (.DIODE(_00475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10379__A2 (.DIODE(_00734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10380__A (.DIODE(_00486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10380__B (.DIODE(_01211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10401__A (.DIODE(_05445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10401__B (.DIODE(_05467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10402__A1 (.DIODE(_05445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10402__A2 (.DIODE(_01177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10402__B2 (.DIODE(_05467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10403__A1 (.DIODE(_01178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10404__A (.DIODE(_02007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10404__B (.DIODE(_02117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10406__A1 (.DIODE(_02029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10406__A2 (.DIODE(_01564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10407__A (.DIODE(_02029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10407__B (.DIODE(_01960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10418__A (.DIODE(_01295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10418__B (.DIODE(_01306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10418__C (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__10419__A1 (.DIODE(_01295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10419__A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__10419__B1 (.DIODE(_02133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10419__B2 (.DIODE(_01306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10420__A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__10421__A (.DIODE(_02127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10421__B (.DIODE(_02459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10423__A1 (.DIODE(_00311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10423__A2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__10424__A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__10425__A (.DIODE(_00322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10425__B (.DIODE(_02673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10452__C (.DIODE(_02703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10453__B1 (.DIODE(_02703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10454__A (.DIODE(_02482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10467__A (.DIODE(_02169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10468__A (.DIODE(_02720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10469__A (.DIODE(_02721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10471__A (.DIODE(_02723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10472__A (.DIODE(_02724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10473__A (.DIODE(_02725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10474__A (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__10475__A (.DIODE(_02727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10476__A (.DIODE(_02728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10477__A (.DIODE(_02730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10478__A1 (.DIODE(_01472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10478__A2 (.DIODE(_02726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10478__B1 (.DIODE(_02731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10478__B2 (.DIODE(_00636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10479__A (.DIODE(_01472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10479__B (.DIODE(_00636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10479__C (.DIODE(_02726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10479__D (.DIODE(_02730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10480__A1 (.DIODE(_02247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10480__A2 (.DIODE(_02722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10481__A (.DIODE(_02726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10482__A (.DIODE(_02735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10483__A (.DIODE(_02731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10484__A (.DIODE(_01473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10484__B (.DIODE(_02247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10484__C (.DIODE(_02736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10484__D (.DIODE(_02737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10485__A1 (.DIODE(_02247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10485__A2 (.DIODE(_02736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10485__B1 (.DIODE(_02737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10485__B2 (.DIODE(_01473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10487__A (.DIODE(_02737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10488__A (.DIODE(_02736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10489__A (.DIODE(_01473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10489__B (.DIODE(_02743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10490__A (.DIODE(_02247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10490__B (.DIODE(_02742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10493__A (.DIODE(_02247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10493__B (.DIODE(_02721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10495__A1 (.DIODE(_00636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10495__A2 (.DIODE(_02735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10495__B1 (.DIODE(_02731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10495__B2 (.DIODE(_00526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10496__A (.DIODE(_00636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10496__B (.DIODE(_00526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10496__C (.DIODE(_02735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10496__D (.DIODE(_02731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10497__A1 (.DIODE(_01473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10497__A2 (.DIODE(_02721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10502__A (.DIODE(_01934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10503__A (.DIODE(_02758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10504__B (.DIODE(_07040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10504__C (.DIODE(_02720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10504__D (.DIODE(_02726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10506__A1 (.DIODE(_00636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10506__A2 (.DIODE(_02721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10506__B1 (.DIODE(_02726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10506__B2 (.DIODE(_00526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10507__A (.DIODE(_01472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10507__B (.DIODE(_02759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10508__A (.DIODE(_02759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10509__A (.DIODE(_02765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10510__A1 (.DIODE(_01473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10510__A2 (.DIODE(_02766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10512__A (.DIODE(_00636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10512__B (.DIODE(_01156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10512__C (.DIODE(_02765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10512__D (.DIODE(_02722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10514__A (.DIODE(_02247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10514__B (.DIODE(_02765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10518__A (.DIODE(_01473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10518__B (.DIODE(_02722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10537__A (.DIODE(_03004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10537__B (.DIODE(_00293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10537__C (.DIODE(_02724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10537__D (.DIODE(_02728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10538__A1 (.DIODE(_00293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10538__A2 (.DIODE(_02725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10538__B1 (.DIODE(_02728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10538__B2 (.DIODE(_03015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10540__A (.DIODE(_00294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10540__B (.DIODE(_02169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10542__A1 (.DIODE(_03004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10542__A2 (.DIODE(_02724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10542__B1 (.DIODE(_02728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10542__B2 (.DIODE(_00388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10543__A (.DIODE(_00388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10543__B (.DIODE(_03004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10543__C (.DIODE(_02724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10543__D (.DIODE(_02727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10544__A1 (.DIODE(_00819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10544__A2 (.DIODE(_02169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10546__A1 (.DIODE(_00818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10546__A2 (.DIODE(_02169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10547__A (.DIODE(_00819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10547__B (.DIODE(_00818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10547__C (.DIODE(_02725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10547__D (.DIODE(_02730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10548__A1 (.DIODE(_00818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10548__A2 (.DIODE(_02725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10548__B1 (.DIODE(_02730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10548__B2 (.DIODE(_00819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10553__A (.DIODE(_00377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10553__B (.DIODE(_02993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10553__C (.DIODE(_02168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10553__D (.DIODE(_02723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10554__A1 (.DIODE(_02993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10554__A2 (.DIODE(_02168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10554__B1 (.DIODE(_02723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10554__B2 (.DIODE(_00377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10555__C (.DIODE(_00095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10555__D (.DIODE(_01933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10558__A (.DIODE(_00293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10558__B (.DIODE(_02169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10560__A (.DIODE(_00294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10560__B (.DIODE(_01934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10564__A1 (.DIODE(_00818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10564__A2 (.DIODE(_02758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10569__A1 (.DIODE(_00819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10569__A2 (.DIODE(_01934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10571__A (.DIODE(_00399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10571__B (.DIODE(_03015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10571__C (.DIODE(_01934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10571__D (.DIODE(_02169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10579__A (.DIODE(_00143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10579__B (.DIODE(_04906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10579__C (.DIODE(_02306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10579__D (.DIODE(_02305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10580__A1 (.DIODE(_00143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10580__A2 (.DIODE(_02306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10580__B1 (.DIODE(_02305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10580__B2 (.DIODE(_04906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10582__A (.DIODE(_00310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10582__B (.DIODE(_01413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10584__A1 (.DIODE(_04895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10584__A2 (.DIODE(_02306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10584__B1 (.DIODE(_02305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10584__B2 (.DIODE(_04928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10585__A (.DIODE(_02158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10586__A (.DIODE(_04895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10586__B (.DIODE(_04928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10586__C (.DIODE(_02849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10586__D (.DIODE(_02304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10587__A1 (.DIODE(_00145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10587__A2 (.DIODE(_01413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10589__A1 (.DIODE(_00310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10589__A2 (.DIODE(_01413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10590__A (.DIODE(_02306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10591__A (.DIODE(_02855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10592__A (.DIODE(_02305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10593__A (.DIODE(_02857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10594__A (.DIODE(_00145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10594__B (.DIODE(_00310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10594__C (.DIODE(_02856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10594__D (.DIODE(_02858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10595__A1 (.DIODE(_00310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10595__A2 (.DIODE(_02855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10595__B1 (.DIODE(_02857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10595__B2 (.DIODE(_00145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10600__A (.DIODE(_04862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10600__B (.DIODE(_04873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10600__C (.DIODE(_01410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10600__D (.DIODE(_02158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10601__A1 (.DIODE(_04862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10601__A2 (.DIODE(_01410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10601__B1 (.DIODE(_02158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10601__B2 (.DIODE(_04873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10602__C (.DIODE(_00142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10602__D (.DIODE(_01059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10605__A (.DIODE(_00144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10605__B (.DIODE(_01412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10607__A (.DIODE(_00158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10607__B (.DIODE(_01059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10611__A1 (.DIODE(_00310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10611__A2 (.DIODE(_01060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10616__A1 (.DIODE(_01472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10616__A2 (.DIODE(_01060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10618__B (.DIODE(_04939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10618__C (.DIODE(_01060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10618__D (.DIODE(_01413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10629__A (.DIODE(_00819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10629__B (.DIODE(_02735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10630__A (.DIODE(_00818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10630__B (.DIODE(_02731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10637__A (.DIODE(_01472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10637__B (.DIODE(_02856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10638__A (.DIODE(_00859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10638__B (.DIODE(_02858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10657__A1 (.DIODE(_00636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10657__A2 (.DIODE(_02765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10657__B1 (.DIODE(_02722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10657__B2 (.DIODE(_01156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10666__A (.DIODE(_00819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10666__B (.DIODE(_00818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10666__C (.DIODE(_02856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10666__D (.DIODE(_02858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10667__A1 (.DIODE(_05192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10667__B2 (.DIODE(_02982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10668__A (.DIODE(_02982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10668__B (.DIODE(_05192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10669__A1 (.DIODE(_05181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10669__A2 (.DIODE(_01411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10670__A (.DIODE(_00094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10670__B (.DIODE(_00151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10670__C (.DIODE(_02849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10670__D (.DIODE(_02304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10671__A1 (.DIODE(_05181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10671__A2 (.DIODE(_02849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10671__B1 (.DIODE(_02304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10671__B2 (.DIODE(_00094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10673__A (.DIODE(_00293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10673__B (.DIODE(_02855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10674__A (.DIODE(_00294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10674__B (.DIODE(_02857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10677__A (.DIODE(_05181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10677__B (.DIODE(_01411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10679__A1 (.DIODE(_02982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10679__B2 (.DIODE(_00377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10680__A (.DIODE(_00366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10680__B (.DIODE(_02982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10681__A1 (.DIODE(_00094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10681__A2 (.DIODE(_01411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10686__A (.DIODE(_05181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10687__A1 (.DIODE(_02982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10687__A2 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__10687__B1 (.DIODE(_02158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10687__B2 (.DIODE(_00366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10688__A (.DIODE(_00366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10688__B (.DIODE(_02982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10688__C (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__10689__A1 (.DIODE(_05203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10692__A (.DIODE(_00094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10692__B (.DIODE(_01411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10701__A (.DIODE(_00095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10701__B (.DIODE(_01059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10703__A (.DIODE(_00388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10703__B (.DIODE(_03004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10703__C (.DIODE(_01059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10703__D (.DIODE(_01412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10722__A1 (.DIODE(_01156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10722__A2 (.DIODE(_02766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10737__A (.DIODE(_00399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10737__B (.DIODE(_03015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10737__C (.DIODE(_02758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10737__D (.DIODE(_02721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10738__A1 (.DIODE(_03015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10738__A2 (.DIODE(_02758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10738__B1 (.DIODE(_02720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10738__B2 (.DIODE(_00399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10742__A2 (.DIODE(_01061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10742__B1 (.DIODE(_01414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10742__B2 (.DIODE(_07040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10753__A1 (.DIODE(_00399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10753__A2 (.DIODE(_02765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10754__A (.DIODE(_00399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10754__B (.DIODE(_02759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10755__A1 (.DIODE(_00526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10755__A2 (.DIODE(_01061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10764__B1 (.DIODE(_01156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10764__C1 (.DIODE(_02766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10765__A1 (.DIODE(_01156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10765__A2 (.DIODE(_02766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10771__B (.DIODE(_06461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10771__C (.DIODE(_02724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10771__D (.DIODE(_02727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10772__A1 (.DIODE(_06461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10772__A2 (.DIODE(_02724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10772__B1 (.DIODE(_02727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10774__A (.DIODE(_06494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10774__B (.DIODE(_02168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10776__A2 (.DIODE(_02723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10776__B1 (.DIODE(_02727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10776__B2 (.DIODE(_02116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10777__A (.DIODE(_02116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10777__B (.DIODE(_02149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10777__C (.DIODE(_02723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10777__D (.DIODE(_02727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10778__A1 (.DIODE(_06937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10778__A2 (.DIODE(_02169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10780__A1 (.DIODE(_06637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10780__A2 (.DIODE(_02720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10781__A (.DIODE(_06937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10781__B (.DIODE(_06494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10781__C (.DIODE(_02725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10781__D (.DIODE(_02730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10782__A1 (.DIODE(_06637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10782__A2 (.DIODE(_02726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10782__B1 (.DIODE(_02730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10782__B2 (.DIODE(_06937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10789__A (.DIODE(_00628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10789__B (.DIODE(_00650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10789__C (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__10791__A1 (.DIODE(_02149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10791__A2 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__10791__B2 (.DIODE(_02105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10792__A (.DIODE(_05588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10792__B (.DIODE(_01933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10793__A1 (.DIODE(_06937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10793__A2 (.DIODE(_02758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10795__A (.DIODE(_02259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10795__B (.DIODE(_02171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10795__C (.DIODE(_02758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10795__D (.DIODE(_02169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10798__A (.DIODE(_06461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10798__B (.DIODE(_02168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10801__A (.DIODE(_06483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10801__B (.DIODE(_01933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10808__A1 (.DIODE(_06494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10808__A2 (.DIODE(_01934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10815__A (.DIODE(_06937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10815__B (.DIODE(_02735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10816__A (.DIODE(_06637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10816__B (.DIODE(_02731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10821__A1 (.DIODE(_00891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10821__A2 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__10821__B1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__10821__B2 (.DIODE(_00989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10822__A (.DIODE(_03587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10822__B (.DIODE(_00891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10822__C (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__10822__D (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__10823__A1 (.DIODE(_01339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10823__A2 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__10824__A (.DIODE(_01372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10824__B (.DIODE(_04268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10824__D (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__10825__A1 (.DIODE(_01339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10825__B1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__10825__B2 (.DIODE(_04081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10828__A (.DIODE(_01383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10828__B (.DIODE(_02724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10829__A (.DIODE(_01350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10829__B (.DIODE(_02728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10830__A1 (.DIODE(_04081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10830__A2 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__10830__B2 (.DIODE(_02727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10832__A (.DIODE(_01339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10832__B (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__10836__A (.DIODE(_01339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10836__B (.DIODE(_01933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10848__A1 (.DIODE(_00541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10848__B1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__10848__B2 (.DIODE(_05742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10849__A (.DIODE(_05742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10849__B (.DIODE(_00541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10849__D (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__10850__A1 (.DIODE(_05566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10850__A2 (.DIODE(_01410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10851__A (.DIODE(_02664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10851__B (.DIODE(_03268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10852__A1 (.DIODE(_03268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10852__A2 (.DIODE(_02158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10852__B1 (.DIODE(_02304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10852__B2 (.DIODE(_05577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10855__A (.DIODE(_06461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10855__B (.DIODE(_02855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10856__A (.DIODE(_06483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10856__B (.DIODE(_02857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10857__A1 (.DIODE(_05588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10857__A2 (.DIODE(_01410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10857__B2 (.DIODE(_02304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10859__A (.DIODE(_03268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10859__B (.DIODE(_01410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10863__A (.DIODE(_05566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10919__A1 (.DIODE(_02171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10919__A2 (.DIODE(_02758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10919__B1 (.DIODE(_02720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10919__B2 (.DIODE(_02467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10926__A (.DIODE(_02467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10926__B (.DIODE(_02758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10950__A (.DIODE(_00143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10950__B (.DIODE(_04906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10950__C (.DIODE(_01508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10950__D (.DIODE(_01504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10951__A1 (.DIODE(_00143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10951__A2 (.DIODE(_01508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10951__B1 (.DIODE(_01505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10951__B2 (.DIODE(_04906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10953__A (.DIODE(_00298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10953__B (.DIODE(_00608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10955__A1 (.DIODE(_04895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10955__A2 (.DIODE(_01507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10955__B1 (.DIODE(_01504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10955__B2 (.DIODE(_04928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10956__A (.DIODE(_04895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10956__B (.DIODE(_04873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10956__C (.DIODE(_01507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10956__D (.DIODE(_01504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10957__A1 (.DIODE(_00145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10957__A2 (.DIODE(_00608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10959__A1 (.DIODE(_00859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10959__A2 (.DIODE(_01400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10960__A (.DIODE(_00145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10960__B (.DIODE(_00310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10960__C (.DIODE(_02187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10960__D (.DIODE(_02189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10961__A1 (.DIODE(_00859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10961__A2 (.DIODE(_02188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10961__B1 (.DIODE(_02190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10961__B2 (.DIODE(_01472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10968__A (.DIODE(_04862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10968__B (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__10968__C (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__10968__D (.DIODE(_01368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10970__A1 (.DIODE(_04862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10970__A2 (.DIODE(_00604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10970__B2 (.DIODE(_04873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10971__A (.DIODE(_00142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10971__B (.DIODE(_00457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10972__A1 (.DIODE(_00145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10972__A2 (.DIODE(_00460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10974__A (.DIODE(_04917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10974__B (.DIODE(_04939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10974__C (.DIODE(_00460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10974__D (.DIODE(_01400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10977__A (.DIODE(_00143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10977__B (.DIODE(_00607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10980__A (.DIODE(_00158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10980__B (.DIODE(_00457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10987__A1 (.DIODE(_00310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10987__A2 (.DIODE(_00459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10994__A (.DIODE(_01473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10994__B (.DIODE(_02188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10995__A (.DIODE(_02247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10995__B (.DIODE(_02190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11000__A1 (.DIODE(_04378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11000__A2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__11000__B1 (.DIODE(_00959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11000__B2 (.DIODE(_02971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11001__A (.DIODE(_02971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11001__B (.DIODE(_04378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11001__C (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__11001__D (.DIODE(_00959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11002__A1 (.DIODE(_05181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11002__A2 (.DIODE(_00604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11003__A (.DIODE(_05192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11003__B (.DIODE(_04598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11003__C (.DIODE(_01368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11003__D (.DIODE(_00959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11004__A1 (.DIODE(_04598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11004__B1 (.DIODE(_01369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11004__B2 (.DIODE(_05203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11007__A (.DIODE(_00293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11007__B (.DIODE(_01664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11008__A (.DIODE(_00294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11008__B (.DIODE(_01505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11009__A1 (.DIODE(_05203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11009__A2 (.DIODE(_00604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11009__B2 (.DIODE(_01369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11011__A (.DIODE(_04598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11011__B (.DIODE(_00604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11015__A (.DIODE(_05181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11015__B (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__11027__A1 (.DIODE(_05027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11027__B2 (.DIODE(_04851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11028__A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__11028__B (.DIODE(_04851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11029__A1 (.DIODE(_00158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11029__A2 (.DIODE(_04037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11030__A (.DIODE(_05027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11030__B (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__11030__C (.DIODE(_00612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11030__D (.DIODE(_00613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11031__A1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__11031__A2 (.DIODE(_00782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11031__B1 (.DIODE(_00778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11031__B2 (.DIODE(_05027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11034__A (.DIODE(_00143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11034__B (.DIODE(_01518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11035__A (.DIODE(_00298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11035__B (.DIODE(_01517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11036__A1 (.DIODE(_00142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11036__A2 (.DIODE(_04037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11036__B2 (.DIODE(_00778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11038__A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__11038__B (.DIODE(_00373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11042__A (.DIODE(_00158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11042__B (.DIODE(_04059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11098__A (.DIODE(_01400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11099__A2 (.DIODE(_01066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11099__B1 (.DIODE(_03414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11099__B2 (.DIODE(_07040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11106__A (.DIODE(_07040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11106__B (.DIODE(_01066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11131__B (.DIODE(_03449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11142__B (.DIODE(_03449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11159__B (.DIODE(_03480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11180__B (.DIODE(_03501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11180__D (.DIODE(_03503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11181__B (.DIODE(_03480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11191__B1 (.DIODE(_01156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11191__C1 (.DIODE(_01108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11192__A1 (.DIODE(_01156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11192__A2 (.DIODE(_01108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11202__B (.DIODE(_03527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11203__B1 (.DIODE(_03503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11203__B2 (.DIODE(_03501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11211__B1 (.DIODE(_02582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11214__B (.DIODE(_03540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11215__B (.DIODE(_03540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11219__A (.DIODE(_00410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11219__B (.DIODE(_01108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11231__B (.DIODE(_03559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11232__B (.DIODE(_03559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11235__A1 (.DIODE(_03015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11235__A2 (.DIODE(_01062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11235__B1 (.DIODE(_01415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11235__B2 (.DIODE(_00410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11237__B (.DIODE(_03566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11242__B (.DIODE(_03571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11249__A (.DIODE(_03566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11259__B (.DIODE(_03571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11260__B (.DIODE(_03527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11296__A (.DIODE(_00819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11296__B (.DIODE(_00818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11296__C (.DIODE(_02736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11296__D (.DIODE(_02737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11339__A (.DIODE(_02673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11340__A (.DIODE(_03678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11341__A (.DIODE(_03679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11342__A (.DIODE(_02459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11343__A (.DIODE(_03681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11344__A (.DIODE(_03682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11345__A (.DIODE(_03683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11346__A (.DIODE(_02135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11347__A (.DIODE(_03686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11348__A1 (.DIODE(_02249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11348__A2 (.DIODE(_01956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11348__B1 (.DIODE(_03687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11348__B2 (.DIODE(_01312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11349__A (.DIODE(_02249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11349__B (.DIODE(_01312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11349__C (.DIODE(_01956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11350__A (.DIODE(_03687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11351__A1 (.DIODE(_00544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11351__B2 (.DIODE(_03690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11352__A (.DIODE(_01155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11352__B (.DIODE(_03680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11353__A (.DIODE(_02246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11353__B (.DIODE(_02249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11353__C (.DIODE(_01956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11353__D (.DIODE(_03687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11354__A1 (.DIODE(_02246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11354__A2 (.DIODE(_01957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11354__B1 (.DIODE(_03690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11354__B2 (.DIODE(_02249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11355__C (.DIODE(_01312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11357__A1_N (.DIODE(_01312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11358__A (.DIODE(_03680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11359__A1 (.DIODE(_01155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11361__A (.DIODE(_00843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11361__B (.DIODE(_00844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11361__C (.DIODE(_03687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11362__A1 (.DIODE(_02246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11362__A2 (.DIODE(_03687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11362__B2 (.DIODE(_02249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11364__A (.DIODE(_01312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11364__B (.DIODE(_03680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11371__A1 (.DIODE(_03690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11372__A (.DIODE(_01155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11374__A (.DIODE(_01312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11374__B (.DIODE(_00544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11374__C (.DIODE(_01957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11374__D (.DIODE(_03690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11381__A1 (.DIODE(_01312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11382__A (.DIODE(_02246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11382__B (.DIODE(_02249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11383__A1 (.DIODE(_02246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11383__B2 (.DIODE(_02249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11392__A (.DIODE(_00112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11392__B (.DIODE(_00268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11392__C (.DIODE(_01179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11392__D (.DIODE(_01254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11393__A1 (.DIODE(_00113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11393__A2 (.DIODE(_01179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11393__B1 (.DIODE(_01249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11393__B2 (.DIODE(_00114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11394__A (.DIODE(_02119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11395__C (.DIODE(_06765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11396__A (.DIODE(_00112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11396__B (.DIODE(_00268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11396__C (.DIODE(_01254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11396__D (.DIODE(_02119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11397__A1 (.DIODE(_00112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11397__A2 (.DIODE(_01254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11397__B1 (.DIODE(_02119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11397__B2 (.DIODE(_00268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11399__A (.DIODE(_02120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11400__A (.DIODE(_00003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11404__A1 (.DIODE(_00004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11404__A2 (.DIODE(_03748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11405__A (.DIODE(_02119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11406__A (.DIODE(_00257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11406__B (.DIODE(_00670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11406__C (.DIODE(_03750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11406__D (.DIODE(_03748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11407__A1 (.DIODE(_00257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11407__A2 (.DIODE(_03750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11407__B1 (.DIODE(_03748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11407__B2 (.DIODE(_00670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11412__A (.DIODE(_00114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11412__B (.DIODE(_06765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11412__C (.DIODE(_01179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11412__D (.DIODE(_01254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11413__A1 (.DIODE(_00268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11413__A2 (.DIODE(_01178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11413__B1 (.DIODE(_01248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11413__B2 (.DIODE(_06733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11415__A (.DIODE(_06775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11415__B (.DIODE(_02119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11417__A1_N (.DIODE(_00003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11419__A (.DIODE(_06775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11422__A1 (.DIODE(_07004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11422__A2 (.DIODE(_03748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11427__A (.DIODE(_00004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11427__B (.DIODE(_06885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11427__C (.DIODE(_01180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11427__D (.DIODE(_01249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11435__A (.DIODE(_03748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11436__A (.DIODE(_03750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11437__A (.DIODE(_00844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11437__B (.DIODE(_03785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11438__A (.DIODE(_00843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11438__B (.DIODE(_03783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11442__A1 (.DIODE(_06964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11442__A2 (.DIODE(_02133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11442__B1 (.DIODE(_02459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11442__B2 (.DIODE(_00121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11443__A (.DIODE(_06964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11443__B (.DIODE(_00121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11443__C (.DIODE(_02133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11443__D (.DIODE(_02459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11444__A1 (.DIODE(_03554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11444__A2 (.DIODE(_03678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11445__A (.DIODE(_00262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11445__B (.DIODE(_00263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11445__C (.DIODE(_03682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11445__D (.DIODE(_03679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11446__A1 (.DIODE(_00262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11446__A2 (.DIODE(_03682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11446__B1 (.DIODE(_03678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11446__B2 (.DIODE(_00263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11448__A (.DIODE(_00263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11448__B (.DIODE(_03683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11449__A (.DIODE(_00262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11449__B (.DIODE(_03680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11451__A (.DIODE(_06964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11451__B (.DIODE(_00121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11451__C (.DIODE(_01953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11451__D (.DIODE(_02133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11452__A1 (.DIODE(_06964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11452__A2 (.DIODE(_01953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11452__B1 (.DIODE(_02134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11452__B2 (.DIODE(_06966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11453__C (.DIODE(_03532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11453__D (.DIODE(_03681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11455__A (.DIODE(_03543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11455__B (.DIODE(_02673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11461__A (.DIODE(_03532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11461__B (.DIODE(_00121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11461__C (.DIODE(_01953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11461__D (.DIODE(_02134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11462__A1 (.DIODE(_00121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11462__A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__11462__B1 (.DIODE(_02133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11462__B2 (.DIODE(_03521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11464__A (.DIODE(_00497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11464__B (.DIODE(_03681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11466__A1_N (.DIODE(_03543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11466__A2_N (.DIODE(_03681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11468__A (.DIODE(_00497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11468__B (.DIODE(_02673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11471__A1 (.DIODE(_00519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11471__A2 (.DIODE(_03679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11476__A (.DIODE(_03554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11476__B (.DIODE(_00508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11476__C (.DIODE(_01954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11476__D (.DIODE(_02135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11527__A1 (.DIODE(_01312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11527__A2 (.DIODE(_01957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11527__B1 (.DIODE(_03690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11527__B2 (.DIODE(_01155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11536__A (.DIODE(_06819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11536__B (.DIODE(_06874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11536__C (.DIODE(_01177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11537__A1 (.DIODE(_06873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11537__A2 (.DIODE(_01178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11537__B2 (.DIODE(_06874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11538__C (.DIODE(_03510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11538__D (.DIODE(_01564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11540__A (.DIODE(_06819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11540__B (.DIODE(_06874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11540__D (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__11541__A1 (.DIODE(_06873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11541__B1 (.DIODE(_01564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11541__B2 (.DIODE(_06874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11543__A (.DIODE(_03521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11543__B (.DIODE(_01960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11546__A1 (.DIODE(_03532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11546__A2 (.DIODE(_02120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11547__A (.DIODE(_06965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11547__B (.DIODE(_06966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11547__C (.DIODE(_02119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11547__D (.DIODE(_02120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11548__A1 (.DIODE(_06964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11548__A2 (.DIODE(_02119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11548__B1 (.DIODE(_02120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11548__B2 (.DIODE(_00121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11553__A1 (.DIODE(_06874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11553__A2 (.DIODE(_01177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11553__B2 (.DIODE(_03510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11554__A (.DIODE(_03510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11554__B (.DIODE(_06874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11554__C (.DIODE(_01177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11555__A1 (.DIODE(_00486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11555__A2 (.DIODE(_01564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11556__A (.DIODE(_00497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11556__B (.DIODE(_02120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11557__A1_N (.DIODE(_03521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11557__A2_N (.DIODE(_02117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11559__A (.DIODE(_00486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11559__B (.DIODE(_01960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11565__A (.DIODE(_00486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11565__B (.DIODE(_02117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11567__A (.DIODE(_03532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11567__B (.DIODE(_00497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11567__C (.DIODE(_01179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11567__D (.DIODE(_01254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11575__A (.DIODE(_00263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11575__B (.DIODE(_03750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11576__A (.DIODE(_00262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11576__B (.DIODE(_03748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11589__A1 (.DIODE(_01155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11589__A2 (.DIODE(_01957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11609__A1 (.DIODE(_00654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11609__A2 (.DIODE(_01181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11609__B1 (.DIODE(_01250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11609__B2 (.DIODE(_00543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11612__A1 (.DIODE(_03554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11612__A2 (.DIODE(_01956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11612__B1 (.DIODE(_03687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11612__B2 (.DIODE(_00519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11620__A1 (.DIODE(_00544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11620__A2 (.DIODE(_01182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11621__A (.DIODE(_00544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11621__B (.DIODE(_01182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11622__A1 (.DIODE(_00519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11622__A2 (.DIODE(_01957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11630__B1 (.DIODE(_01155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11630__C1 (.DIODE(_01958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11631__A1 (.DIODE(_01155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11631__A2 (.DIODE(_01957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11646__A (.DIODE(_02249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11647__A (.DIODE(_02246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11662__A (.DIODE(_00258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11662__B (.DIODE(_06765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11662__C (.DIODE(_00414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11663__A1 (.DIODE(_00258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11663__A2 (.DIODE(_00414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11663__B1 (.DIODE(_00574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11663__B2 (.DIODE(_06765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11664__A1 (.DIODE(_00575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11665__A (.DIODE(_06885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11665__B (.DIODE(_01601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11667__A (.DIODE(_00004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11667__B (.DIODE(_06885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11667__C (.DIODE(_00416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11667__D (.DIODE(_01288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11669__A1 (.DIODE(_06733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11669__A2 (.DIODE(_03773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11669__B2 (.DIODE(_03696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11670__A (.DIODE(_07010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11670__B (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__11670__C (.DIODE(_03718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11670__D (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__11671__A1 (.DIODE(_07010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11671__A2 (.DIODE(_00423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11671__B1 (.DIODE(_03762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11671__B2 (.DIODE(_00101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11672__C (.DIODE(_06733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11672__D (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__11673__A1_N (.DIODE(_06733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11673__A2_N (.DIODE(_03938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11676__A (.DIODE(_00112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11676__B (.DIODE(_00268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11676__C (.DIODE(_00755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11676__D (.DIODE(_01260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11677__A1 (.DIODE(_07010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11677__A2 (.DIODE(_03773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11677__B1 (.DIODE(_01260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11677__B2 (.DIODE(_00268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11688__A1 (.DIODE(_03510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11688__A2 (.DIODE(_00734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11688__B2 (.DIODE(_00413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11689__A (.DIODE(_06819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11689__B (.DIODE(_06821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11689__C (.DIODE(_00730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11689__D (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__11690__A1 (.DIODE(_06819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11690__A2 (.DIODE(_00571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11690__B1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__11690__B2 (.DIODE(_06874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11691__C (.DIODE(_03510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11691__D (.DIODE(_01211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11692__A1_N (.DIODE(_03510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11692__A2_N (.DIODE(_01211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11695__A (.DIODE(_06964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11695__B (.DIODE(_06875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11695__C (.DIODE(_01272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11695__D (.DIODE(_01211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11696__A1 (.DIODE(_06873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11696__A2 (.DIODE(_01272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11696__B1 (.DIODE(_01211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11696__B2 (.DIODE(_06875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11710__A (.DIODE(_00258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11710__B (.DIODE(_00915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11711__A (.DIODE(_00257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11711__B (.DIODE(_00916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11718__A (.DIODE(_00263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11718__B (.DIODE(_01600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11719__A (.DIODE(_00262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11719__B (.DIODE(_01585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11739__A1 (.DIODE(_00654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11739__A2 (.DIODE(_01188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11739__B1 (.DIODE(_01289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11739__B2 (.DIODE(_00543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11746__A (.DIODE(_00543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11746__B (.DIODE(_01188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11762__A (.DIODE(_00138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11762__B (.DIODE(_02018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11762__C (.DIODE(_01953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11763__A1 (.DIODE(_00138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11763__A2 (.DIODE(_01953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11763__B1 (.DIODE(_02134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11763__B2 (.DIODE(_02018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11764__A1 (.DIODE(_02135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11765__A (.DIODE(_02280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11765__B (.DIODE(_03682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11767__A (.DIODE(_03070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11767__B (.DIODE(_02335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11767__C (.DIODE(_01954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11767__D (.DIODE(_02135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11769__A1 (.DIODE(_02007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11769__A2 (.DIODE(_01564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11769__B2 (.DIODE(_01178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11770__A (.DIODE(_05445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11770__B (.DIODE(_05731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11770__D (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__11771__A1 (.DIODE(_05445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11771__B1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__11771__B2 (.DIODE(_05467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11772__C (.DIODE(_01996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11772__D (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__11773__A1_N (.DIODE(_01996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11773__A2_N (.DIODE(_01960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11776__A (.DIODE(_05456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11776__B (.DIODE(_05478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11776__C (.DIODE(_02117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11776__D (.DIODE(_01960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11777__A1 (.DIODE(_05456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11777__A2 (.DIODE(_02117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11777__B1 (.DIODE(_01960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11777__B2 (.DIODE(_05478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11788__A1 (.DIODE(_02127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11788__A2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__11788__B2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__11789__C (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__11789__D (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__11790__A1 (.DIODE(_01295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11790__A2 (.DIODE(_02133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11790__B1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__11790__B2 (.DIODE(_01306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11791__C (.DIODE(_01744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11791__D (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__11792__A1_N (.DIODE(_02127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11792__A2_N (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__11795__A (.DIODE(_01361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11795__B (.DIODE(_00159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11795__C (.DIODE(_02459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11795__D (.DIODE(_02673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11796__A1 (.DIODE(_01361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11796__A2 (.DIODE(_02459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11796__B1 (.DIODE(_02673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11796__B2 (.DIODE(_01405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11810__A (.DIODE(_06439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11810__B (.DIODE(_03750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11811__A (.DIODE(_06428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11811__B (.DIODE(_03748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11818__A (.DIODE(_00159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11818__B (.DIODE(_03682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11819__A (.DIODE(_00157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11819__B (.DIODE(_03678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11839__A1 (.DIODE(_03070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11839__A2 (.DIODE(_01955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11839__B1 (.DIODE(_03686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11839__B2 (.DIODE(_02456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11846__A (.DIODE(_02456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11846__B (.DIODE(_01955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11866__A (.DIODE(_00113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11866__B (.DIODE(_00258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11866__C (.DIODE(_00415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11866__D (.DIODE(_00574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11867__A1 (.DIODE(_00113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11867__A2 (.DIODE(_00415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11867__B1 (.DIODE(_00575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11867__B2 (.DIODE(_00258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11868__C (.DIODE(_00003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11868__D (.DIODE(_01600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11869__A1 (.DIODE(_06775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11869__A2 (.DIODE(_01600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11869__B2 (.DIODE(_00575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11870__A (.DIODE(_06885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11870__B (.DIODE(_01780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11871__A1_N (.DIODE(_00004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11871__A2_N (.DIODE(_01601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11872__A1 (.DIODE(_07004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11872__A2 (.DIODE(_01780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11880__A (.DIODE(_00257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11880__B (.DIODE(_00670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11880__C (.DIODE(_00915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11880__D (.DIODE(_00916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11882__A (.DIODE(_00262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11882__B (.DIODE(_00263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11882__C (.DIODE(_02090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11882__D (.DIODE(_01780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11897__A (.DIODE(_06417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11897__B (.DIODE(_06439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11897__C (.DIODE(_01954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11897__D (.DIODE(_02135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11898__A1 (.DIODE(_06428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11898__A2 (.DIODE(_01954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11898__B1 (.DIODE(_02135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11898__B2 (.DIODE(_06439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11899__C (.DIODE(_03059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11899__D (.DIODE(_03682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11900__A1 (.DIODE(_02040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11900__A2 (.DIODE(_03681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11900__B2 (.DIODE(_02135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11901__A (.DIODE(_02280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11901__B (.DIODE(_03678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11902__A1_N (.DIODE(_03070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11902__A2_N (.DIODE(_03682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11903__A1 (.DIODE(_02335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11903__A2 (.DIODE(_03678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11911__A (.DIODE(_06626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11911__B (.DIODE(_06450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11911__C (.DIODE(_03750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11911__D (.DIODE(_03783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11913__A (.DIODE(_00157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11913__B (.DIODE(_00159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11913__C (.DIODE(_03683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11913__D (.DIODE(_03679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11931__A (.DIODE(_00113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11931__B (.DIODE(_00114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11931__C (.DIODE(_00572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11931__D (.DIODE(_01272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11932__A (.DIODE(_00114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11932__B (.DIODE(_01272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11933__A1 (.DIODE(_00113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11933__A2 (.DIODE(_00574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11935__A (.DIODE(_00003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11935__B (.DIODE(_01585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11936__A1 (.DIODE(_00004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11936__A2 (.DIODE(_01585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11957__A (.DIODE(_06417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11957__B (.DIODE(_00138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11957__C (.DIODE(_02134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11957__D (.DIODE(_03681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11958__A (.DIODE(_00138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11958__B (.DIODE(_02459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11959__A1 (.DIODE(_06417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11959__A2 (.DIODE(_02134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11961__A (.DIODE(_03059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11961__B (.DIODE(_03678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11962__A1 (.DIODE(_03059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11962__A2 (.DIODE(_03678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11990__B1 (.DIODE(_00530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11990__C1 (.DIODE(_01958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11991__A1 (.DIODE(_00530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11991__A2 (.DIODE(_01958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12004__A (.DIODE(_00257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12004__B (.DIODE(_00670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12004__C (.DIODE(_02090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12004__D (.DIODE(_01780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12005__A1 (.DIODE(_00843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12005__A2 (.DIODE(_02090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12005__B1 (.DIODE(_02088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12005__B2 (.DIODE(_00844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12022__A (.DIODE(_06626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12022__B (.DIODE(_06450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12022__C (.DIODE(_03683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12022__D (.DIODE(_03679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12023__A1 (.DIODE(_06626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12023__A2 (.DIODE(_03683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12023__B1 (.DIODE(_03679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12023__B2 (.DIODE(_06450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12068__A1 (.DIODE(_03554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12068__A2 (.DIODE(_01183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12068__B1 (.DIODE(_01252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12068__B2 (.DIODE(_00530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12080__A (.DIODE(_02246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12080__B (.DIODE(_02426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12090__A (.DIODE(_06626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12090__B (.DIODE(_03680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12144__A (.DIODE(_00530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12144__B (.DIODE(_01183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12178__B (.DIODE(_04600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12203__B (.DIODE(_04627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12205__A (.DIODE(_00374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12205__B (.DIODE(_00784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12205__C (.DIODE(_01953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12205__D (.DIODE(_02134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12206__A1 (.DIODE(_00784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12206__A2 (.DIODE(_01953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12206__B1 (.DIODE(_02134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12206__B2 (.DIODE(_00374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12207__B (.DIODE(_03682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12207__C (.DIODE(_00379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12208__A1 (.DIODE(_01518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12208__A2 (.DIODE(_01954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12208__B1 (.DIODE(_02135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12209__A1_N (.DIODE(_00379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12209__A2_N (.DIODE(_03682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12211__A (.DIODE(_00376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12211__B (.DIODE(_00379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12211__C (.DIODE(_01954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12211__D (.DIODE(_02135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12213__A (.DIODE(_00605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12213__B (.DIODE(_01507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12213__C (.DIODE(_01179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12213__D (.DIODE(_01254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12214__A1 (.DIODE(_01507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12214__A2 (.DIODE(_01179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12214__B1 (.DIODE(_01254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12214__B2 (.DIODE(_00605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12215__B (.DIODE(_03750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12215__C (.DIODE(_00458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12216__A1 (.DIODE(_01664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12216__A2 (.DIODE(_01180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12216__B1 (.DIODE(_01249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12216__B2 (.DIODE(_00607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12217__A1_N (.DIODE(_00458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12217__A2_N (.DIODE(_03750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12219__A (.DIODE(_00459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12219__B (.DIODE(_00608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12219__C (.DIODE(_01180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12219__D (.DIODE(_01249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12223__A1 (.DIODE(_00778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12223__A2 (.DIODE(_01248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12223__B1 (.DIODE(_02117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12223__B2 (.DIODE(_00783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12224__A (.DIODE(_00783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12224__B (.DIODE(_00778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12224__C (.DIODE(_01248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12224__D (.DIODE(_02117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12226__A (.DIODE(_01518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12226__B (.DIODE(_01517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12227__A1 (.DIODE(_01517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12227__B2 (.DIODE(_01518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12229__A (.DIODE(_01518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12229__B (.DIODE(_03750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12230__A (.DIODE(_01517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12230__B (.DIODE(_03748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12234__A1 (.DIODE(_00778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12234__A2 (.DIODE(_01178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12234__B1 (.DIODE(_01248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12234__B2 (.DIODE(_00783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12235__A (.DIODE(_00783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12235__B (.DIODE(_00778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12235__C (.DIODE(_01178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12235__D (.DIODE(_01248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12236__A2 (.DIODE(_03750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12238__B (.DIODE(_02120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12245__A1 (.DIODE(_00783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12245__A2 (.DIODE(_01178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12245__B1 (.DIODE(_01248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12245__B2 (.DIODE(_04037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12246__A (.DIODE(_04037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12246__B (.DIODE(_00783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12246__C (.DIODE(_01178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12246__D (.DIODE(_01248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12247__A1 (.DIODE(_00378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12247__A2 (.DIODE(_02119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12248__A (.DIODE(_00379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12248__B (.DIODE(_03748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12252__A (.DIODE(_00378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12252__B (.DIODE(_02120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12258__A (.DIODE(_00378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12260__A (.DIODE(_00376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12260__B (.DIODE(_00378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12260__C (.DIODE(_01180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12260__D (.DIODE(_01249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12270__A1 (.DIODE(_03414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12270__A2 (.DIODE(_01181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12270__B1 (.DIODE(_01250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12270__B2 (.DIODE(_01066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12274__A1 (.DIODE(_00376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12274__A2 (.DIODE(_01955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12274__B1 (.DIODE(_03686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12274__B2 (.DIODE(_00380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12281__A (.DIODE(_01066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12284__A1 (.DIODE(_04714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12284__A2 (.DIODE(_01182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12285__A (.DIODE(_04714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12285__B (.DIODE(_01181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12286__A1 (.DIODE(_00380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12286__A2 (.DIODE(_01956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12292__A1 (.DIODE(_02187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12292__A2 (.DIODE(_01601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12292__B1 (.DIODE(_02189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12292__B2 (.DIODE(_00575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12293__A (.DIODE(_00575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12293__B (.DIODE(_01664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12293__C (.DIODE(_01601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12293__D (.DIODE(_01505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12294__A1 (.DIODE(_03414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12294__A2 (.DIODE(_02426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12295__A (.DIODE(_02188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12295__B (.DIODE(_02427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12295__C (.DIODE(_02190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12295__D (.DIODE(_02088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12296__A1 (.DIODE(_02427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12296__A2 (.DIODE(_02190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12296__B1 (.DIODE(_02088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12296__B2 (.DIODE(_02188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12299__A (.DIODE(_02188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12299__B (.DIODE(_02427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12300__A (.DIODE(_02190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12300__B (.DIODE(_02426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12302__A (.DIODE(_00415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12302__B (.DIODE(_00575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12302__C (.DIODE(_01664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12302__D (.DIODE(_01505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12303__A1 (.DIODE(_01288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12303__A2 (.DIODE(_02187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12303__B1 (.DIODE(_02189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12303__B2 (.DIODE(_00416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12304__C (.DIODE(_00608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12304__D (.DIODE(_01601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12306__A (.DIODE(_01400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12306__B (.DIODE(_01780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12311__A1 (.DIODE(_00607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12311__A2 (.DIODE(_00575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12311__B1 (.DIODE(_01664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12311__B2 (.DIODE(_00415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12312__A (.DIODE(_00415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12312__B (.DIODE(_00607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12312__C (.DIODE(_01664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12313__A1 (.DIODE(_00459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12313__A2 (.DIODE(_01601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12313__B2 (.DIODE(_01288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12314__A (.DIODE(_00459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12314__B (.DIODE(_01780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12315__A1_N (.DIODE(_00608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12315__A2_N (.DIODE(_01601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12317__A1 (.DIODE(_00460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12317__A2 (.DIODE(_02088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12325__A1 (.DIODE(_01289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12326__A (.DIODE(_00460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12326__B (.DIODE(_02090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12328__A (.DIODE(_01066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12328__B (.DIODE(_01188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12328__C (.DIODE(_03414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12328__D (.DIODE(_01289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12339__A (.DIODE(_00755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12339__B (.DIODE(_01260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12339__C (.DIODE(_01507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12339__D (.DIODE(_01369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12340__A1 (.DIODE(_03762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12340__A2 (.DIODE(_01368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12340__B1 (.DIODE(_00959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12341__B (.DIODE(_03762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12341__C (.DIODE(_01368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12341__D (.DIODE(_00959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12342__A1 (.DIODE(_01260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12342__A2 (.DIODE(_00605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12343__A1 (.DIODE(_01260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12343__B1 (.DIODE(_01369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12343__B2 (.DIODE(_00755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12345__A (.DIODE(_00915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12345__B (.DIODE(_01664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12346__A (.DIODE(_00916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12346__B (.DIODE(_01505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12349__A (.DIODE(_01260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12349__B (.DIODE(_00605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12351__B1 (.DIODE(_01369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12351__B2 (.DIODE(_03696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12352__A (.DIODE(_03696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12352__D (.DIODE(_01369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12353__A1 (.DIODE(_00742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12353__A2 (.DIODE(_00605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12359__A (.DIODE(_00742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12359__B (.DIODE(_00605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12361__A2 (.DIODE(_00604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12361__B2 (.DIODE(_03696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12362__A (.DIODE(_03696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12362__C (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__12363__A1 (.DIODE(_00755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12363__A2 (.DIODE(_00457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12364__A (.DIODE(_00741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12364__B (.DIODE(_00457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12372__A (.DIODE(_00914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12372__B (.DIODE(_00457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12374__A (.DIODE(_00389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12374__B (.DIODE(_00392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12374__C (.DIODE(_00457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12374__D (.DIODE(_00607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12385__A1 (.DIODE(_00778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12385__A2 (.DIODE(_00571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12385__B1 (.DIODE(_00734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12385__B2 (.DIODE(_00782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12386__A (.DIODE(_00782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12386__B (.DIODE(_00613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12386__C (.DIODE(_00571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12386__D (.DIODE(_00734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12387__A1 (.DIODE(_00374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12387__A2 (.DIODE(_01584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12388__A (.DIODE(_00784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12388__B (.DIODE(_00779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12388__C (.DIODE(_01586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12388__D (.DIODE(_01584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12389__A1 (.DIODE(_00779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12389__A2 (.DIODE(_01586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12389__B1 (.DIODE(_01584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12389__B2 (.DIODE(_00784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12391__A (.DIODE(_01518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12391__B (.DIODE(_01601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12392__A (.DIODE(_01517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12392__B (.DIODE(_01780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12394__A1 (.DIODE(_00778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12394__A2 (.DIODE(_00413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12394__B1 (.DIODE(_00571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12394__B2 (.DIODE(_00782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12395__A (.DIODE(_00782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12395__B (.DIODE(_00613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12395__C (.DIODE(_00413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12395__D (.DIODE(_00571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12396__A1 (.DIODE(_00374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12396__A2 (.DIODE(_01272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12398__A (.DIODE(_00374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12398__B (.DIODE(_01584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12404__A (.DIODE(_00374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12404__B (.DIODE(_01272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12406__A1 (.DIODE(_00782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12406__A2 (.DIODE(_00413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12406__B1 (.DIODE(_00571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12406__B2 (.DIODE(_00373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12407__A (.DIODE(_00373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12407__B (.DIODE(_00782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12407__C (.DIODE(_00413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12407__D (.DIODE(_00571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12408__A1 (.DIODE(_04059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12408__A2 (.DIODE(_01272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12409__A (.DIODE(_04059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12409__B (.DIODE(_01584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12411__A (.DIODE(_00378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12411__B (.DIODE(_01584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12416__A (.DIODE(_00378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12416__B (.DIODE(_01586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12418__B (.DIODE(_00378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12418__C (.DIODE(_00414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12418__D (.DIODE(_00572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12470__A1 (.DIODE(_02008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12470__A2 (.DIODE(_03414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12470__B1 (.DIODE(_01289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12470__B2 (.DIODE(_04714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12477__A (.DIODE(_04714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12477__B (.DIODE(_02008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12482__B1 (.DIODE(_03762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12482__B2 (.DIODE(_00612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12483__A (.DIODE(_00612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12483__C (.DIODE(_00423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12483__D (.DIODE(_03762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12484__A1 (.DIODE(_00374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12484__A2 (.DIODE(_00741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12485__A (.DIODE(_00784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12485__B (.DIODE(_00779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12485__C (.DIODE(_00742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12485__D (.DIODE(_00741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12486__A1 (.DIODE(_00779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12486__A2 (.DIODE(_00755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12486__B1 (.DIODE(_00741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12486__B2 (.DIODE(_00783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12488__A (.DIODE(_01518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12488__B (.DIODE(_00914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12489__A (.DIODE(_01517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12489__B (.DIODE(_00916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12491__A1 (.DIODE(_00613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12491__A2 (.DIODE(_03696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12491__B2 (.DIODE(_00612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12492__C (.DIODE(_03685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12492__D (.DIODE(_00423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12493__A1 (.DIODE(_00374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12493__A2 (.DIODE(_00755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12495__A (.DIODE(_04037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12495__B (.DIODE(_03938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12500__A1 (.DIODE(_00612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12500__A2 (.DIODE(_03696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12500__B2 (.DIODE(_04026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12501__A (.DIODE(_04026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12501__C (.DIODE(_03685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12501__D (.DIODE(_00423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12502__A1 (.DIODE(_04048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12502__A2 (.DIODE(_03894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12503__A (.DIODE(_00378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12503__B (.DIODE(_00741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12505__A (.DIODE(_04037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12505__B (.DIODE(_03773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12507__A (.DIODE(_04059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12507__B (.DIODE(_03938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12513__A (.DIODE(_04059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12513__B (.DIODE(_00755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12515__A (.DIODE(_00374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12515__B (.DIODE(_04059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12515__C (.DIODE(_03707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12515__D (.DIODE(_03740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12546__A1 (.DIODE(_00393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12546__A2 (.DIODE(_00459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12546__B1 (.DIODE(_01400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12546__B2 (.DIODE(_00390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12551__A1 (.DIODE(_00376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12551__A2 (.DIODE(_01188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12551__B1 (.DIODE(_01289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12551__B2 (.DIODE(_00380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12560__A1 (.DIODE(_00390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12560__A2 (.DIODE(_04714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12561__A (.DIODE(_00390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12561__B (.DIODE(_01066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12562__A1 (.DIODE(_00380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12562__A2 (.DIODE(_02008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12577__A (.DIODE(_00389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12577__B (.DIODE(_00393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12577__C (.DIODE(_01934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12577__D (.DIODE(_02169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12579__A1 (.DIODE(_00393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12579__A2 (.DIODE(_02758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12579__B1 (.DIODE(_02720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12579__B2 (.DIODE(_00390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12580__A (.DIODE(_03740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12580__B (.DIODE(_00742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12580__C (.DIODE(_02849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12580__D (.DIODE(_02304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12581__A1 (.DIODE(_00742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12581__A2 (.DIODE(_02849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12581__B1 (.DIODE(_02304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12581__B2 (.DIODE(_00392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12583__A (.DIODE(_00745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12583__B (.DIODE(_01412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12585__A1 (.DIODE(_03740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12585__A2 (.DIODE(_02158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12585__B1 (.DIODE(_02304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12585__B2 (.DIODE(_03707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12586__A (.DIODE(_03707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12586__B (.DIODE(_03740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12586__C (.DIODE(_02158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12586__D (.DIODE(_02304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12587__A1 (.DIODE(_00915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12587__A2 (.DIODE(_01412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12589__A1 (.DIODE(_00745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12589__A2 (.DIODE(_01412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12590__A (.DIODE(_00915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12590__B (.DIODE(_00916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12590__C (.DIODE(_02855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12590__D (.DIODE(_02857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12591__A1 (.DIODE(_00745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12591__A2 (.DIODE(_02855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12591__B1 (.DIODE(_02857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12591__B2 (.DIODE(_00914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12596__A (.DIODE(_00745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12596__B (.DIODE(_01059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12597__A1 (.DIODE(_03740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12597__A2 (.DIODE(_01411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12597__B1 (.DIODE(_02849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12597__B2 (.DIODE(_03707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12598__A (.DIODE(_03707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12598__B (.DIODE(_03740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12598__C (.DIODE(_01411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12598__D (.DIODE(_02849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12599__A1 (.DIODE(_00914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12599__A2 (.DIODE(_01059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12602__A (.DIODE(_00914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12602__B (.DIODE(_01412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12609__A (.DIODE(_00915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12609__B (.DIODE(_01059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12611__A (.DIODE(_00389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12611__B (.DIODE(_00393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12611__C (.DIODE(_01060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12611__D (.DIODE(_01412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12619__A (.DIODE(_00415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12619__B (.DIODE(_00575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12619__C (.DIODE(_01060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12619__D (.DIODE(_01413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12620__A1 (.DIODE(_01289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12620__A2 (.DIODE(_01061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12620__B1 (.DIODE(_01414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12620__B2 (.DIODE(_01188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12624__A (.DIODE(_00414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12624__B (.DIODE(_00572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12624__C (.DIODE(_02849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12625__A1 (.DIODE(_00572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12625__A2 (.DIODE(_01411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12625__B1 (.DIODE(_02306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12625__B2 (.DIODE(_00414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12626__A1 (.DIODE(_01413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12627__A (.DIODE(_01600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12627__B (.DIODE(_01060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12632__A (.DIODE(_00389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12632__B (.DIODE(_00392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12632__C (.DIODE(_02723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12633__A1 (.DIODE(_00392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12633__A2 (.DIODE(_02168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12633__B1 (.DIODE(_02723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12633__B2 (.DIODE(_00389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12634__A1 (.DIODE(_02168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12635__A (.DIODE(_00915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12635__B (.DIODE(_01933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12640__A (.DIODE(_00915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12640__B (.DIODE(_02855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12641__A (.DIODE(_00916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12641__B (.DIODE(_02857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12649__A (.DIODE(_02008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12649__B (.DIODE(_01061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12652__A (.DIODE(_00390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12652__B (.DIODE(_02759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12654__A1 (.DIODE(_00390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12654__A2 (.DIODE(_02759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12666__B1_N (.DIODE(_05136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12675__B1 (.DIODE(_00381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12675__C1 (.DIODE(_01958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12676__A1 (.DIODE(_00381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12676__A2 (.DIODE(_01958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12679__A (.DIODE(_05136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12681__A2 (.DIODE(_05150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12684__C (.DIODE(_05150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12685__B1 (.DIODE(_05150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12711__A1 (.DIODE(_00393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12711__A2 (.DIODE(_01062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12711__B1 (.DIODE(_01415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12711__B2 (.DIODE(_00391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12714__A1 (.DIODE(_00376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12714__A2 (.DIODE(_01183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12714__B1 (.DIODE(_01252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12714__B2 (.DIODE(_00380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12719__A (.DIODE(_05193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12721__A (.DIODE(_00391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12721__B (.DIODE(_01108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12722__A (.DIODE(_00380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12722__B (.DIODE(_01182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12723__A1 (.DIODE(_00391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12723__A2 (.DIODE(_01062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12729__A (.DIODE(_05193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12735__A2 (.DIODE(_05150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12741__A (.DIODE(_00783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12741__B (.DIODE(_00779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12741__C (.DIODE(_02133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12742__A1 (.DIODE(_00779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12742__A2 (.DIODE(_01953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12742__B1 (.DIODE(_02134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12742__B2 (.DIODE(_00784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12743__A1 (.DIODE(_01953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12744__B (.DIODE(_03681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12746__A1 (.DIODE(_00378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12746__A2 (.DIODE(_03681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12747__A (.DIODE(_00379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12747__B (.DIODE(_03678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12753__A (.DIODE(_01507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12753__B (.DIODE(_01504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12753__C (.DIODE(_01248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12754__A1 (.DIODE(_01504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12754__A2 (.DIODE(_01179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12754__B1 (.DIODE(_01254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12754__B2 (.DIODE(_01507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12755__A1 (.DIODE(_01180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12756__A (.DIODE(_00607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12758__A1 (.DIODE(_00457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12759__A (.DIODE(_00457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12780__A1 (.DIODE(_00572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12780__A2 (.DIODE(_02849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12780__B1 (.DIODE(_02305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12780__B2 (.DIODE(_00414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12781__A1 (.DIODE(_02305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12782__A (.DIODE(_01600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12782__B (.DIODE(_01412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12784__A (.DIODE(_00414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12784__B (.DIODE(_00572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12784__C (.DIODE(_01411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12784__D (.DIODE(_02849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12785__A1 (.DIODE(_01586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12785__A2 (.DIODE(_01059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12786__A (.DIODE(_01585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12786__B (.DIODE(_01059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12792__A1 (.DIODE(_00392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12792__A2 (.DIODE(_02723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12792__B1 (.DIODE(_02727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12792__B2 (.DIODE(_00389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12793__A1 (.DIODE(_02728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12794__A (.DIODE(_00914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12794__B (.DIODE(_02168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12796__A (.DIODE(_00389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12796__B (.DIODE(_00392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12796__C (.DIODE(_02168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12796__D (.DIODE(_02723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12797__A1 (.DIODE(_00914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12797__A2 (.DIODE(_01933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12798__A (.DIODE(_00916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12798__B (.DIODE(_01933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12830__B1 (.DIODE(_04600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12835__A (.DIODE(_00916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12835__B (.DIODE(_01933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12837__A1_N (.DIODE(_02728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12838__A1 (.DIODE(_00742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12838__A2 (.DIODE(_02724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12838__B1 (.DIODE(_02727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12838__B2 (.DIODE(_00392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12839__A (.DIODE(_00392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12839__B (.DIODE(_00742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12839__C (.DIODE(_02723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12839__D (.DIODE(_02727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12841__A (.DIODE(_00745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12841__B (.DIODE(_02168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12849__A (.DIODE(_01585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12849__B (.DIODE(_01060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12851__A1_N (.DIODE(_02857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12852__A1 (.DIODE(_01586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12852__A2 (.DIODE(_02306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12852__B1 (.DIODE(_02305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12852__B2 (.DIODE(_00574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12853__A (.DIODE(_00572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12853__B (.DIODE(_01586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12853__C (.DIODE(_02306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12853__D (.DIODE(_02305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12855__A (.DIODE(_01584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12855__B (.DIODE(_01412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12866__A (.DIODE(_02008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12866__B (.DIODE(_02765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12873__A (.DIODE(_00458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12873__B (.DIODE(_03748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12875__A1_N (.DIODE(_01180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12876__A (.DIODE(_01504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12876__B (.DIODE(_01249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12877__A (.DIODE(_01507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12877__B (.DIODE(_02119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12878__A (.DIODE(_01507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12878__B (.DIODE(_01369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12878__C (.DIODE(_01248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12878__D (.DIODE(_02117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12880__A (.DIODE(_00605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12880__B (.DIODE(_02120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12888__A (.DIODE(_00379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12888__B (.DIODE(_03678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12890__A1_N (.DIODE(_01954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12891__A (.DIODE(_00779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12891__B (.DIODE(_02134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12892__A (.DIODE(_00784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12892__B (.DIODE(_02459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12893__A (.DIODE(_00783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12893__B (.DIODE(_00778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12893__C (.DIODE(_02133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12893__D (.DIODE(_02459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12895__B (.DIODE(_02673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12908__A (.DIODE(_04714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12908__B (.DIODE(_01957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12918__A (.DIODE(_01108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12918__B (.DIODE(_01183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12932__B (.DIODE(_05429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12942__A2 (.DIODE(_02150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12948__B (.DIODE(_05447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12953__A2 (.DIODE(_05451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12956__B (.DIODE(_05429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12966__A (.DIODE(_05464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12969__A (.DIODE(_05455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12972__A (.DIODE(_05451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12973__B (.DIODE(_05447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12981__B (.DIODE(_05483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12986__A2 (.DIODE(_05487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12991__B (.DIODE(_05483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12992__A2 (.DIODE(_05494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12994__B1 (.DIODE(_00381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12994__C1 (.DIODE(_02008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12995__A1 (.DIODE(_00381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12995__A2 (.DIODE(_02008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12997__A2 (.DIODE(_05494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12997__B1 (.DIODE(_05501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12999__A (.DIODE(_05487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13005__B (.DIODE(_05494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13010__B (.DIODE(_05513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13010__D (.DIODE(_05515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13013__A1 (.DIODE(_05509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13014__B (.DIODE(_05494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13016__A (.DIODE(_05501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13018__B (.DIODE(_05507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13018__C (.DIODE(_05524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13023__A (.DIODE(_05509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13024__B1 (.DIODE(_05515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13024__B2 (.DIODE(_05513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13031__A (.DIODE(_05536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13034__B1 (.DIODE(_05541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13039__A (.DIODE(_05541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13040__A (.DIODE(_05536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13046__B (.DIODE(_05554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13048__A1 (.DIODE(_00376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13048__A2 (.DIODE(_00391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13048__B1 (.DIODE(_00393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13048__B2 (.DIODE(_00381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13050__B1 (.DIODE(_05559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13053__A (.DIODE(_05546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13054__B (.DIODE(_05554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13056__A2 (.DIODE(_02703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13058__A (.DIODE(_00381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13058__B (.DIODE(_00391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13061__A (.DIODE(_05559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13081__B1 (.DIODE(_05593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13090__A2 (.DIODE(_05595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13091__B (.DIODE(_04627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13106__B (.DIODE(_05620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13120__B (.DIODE(_05636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13121__B (.DIODE(_05620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13134__B (.DIODE(_05651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13135__B (.DIODE(_05636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13148__B (.DIODE(_05651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13151__B (.DIODE(_05670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13162__B (.DIODE(_05670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13167__B (.DIODE(_05688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13182__B (.DIODE(_05704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13183__B (.DIODE(_05688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13192__A (.DIODE(_05464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13194__B (.DIODE(_05704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13203__A1 (.DIODE(_05455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13227__A (.DIODE(_05424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13233__A1 (.DIODE(_02278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13251__A (.DIODE(_05776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13251__B (.DIODE(_05773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13252__A (.DIODE(_05546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13253__A (.DIODE(_05524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13255__A (.DIODE(_05524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13255__B (.DIODE(_05546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13256__B (.DIODE(_05779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13260__A2 (.DIODE(_05779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13260__B1 (.DIODE(_05784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13261__A1 (.DIODE(_02278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13262__B (.DIODE(_05786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13264__A (.DIODE(_05507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13264__B (.DIODE(_05524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13265__A1 (.DIODE(_05507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13265__A2 (.DIODE(_05524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13265__A3 (.DIODE(_05593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13266__B1 (.DIODE(_05789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13268__B (.DIODE(_05792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13270__A (.DIODE(_05779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13271__A1 (.DIODE(_05773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13271__A2 (.DIODE(_05776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13274__A1 (.DIODE(_05784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13283__A1 (.DIODE(_05786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13286__B (.DIODE(_05807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13289__A (.DIODE(_05789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13289__B (.DIODE(_05807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13290__A (.DIODE(_05810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13303__A2 (.DIODE(_05595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13311__A1 (.DIODE(_05786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13312__B (.DIODE(_05833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13319__A1 (.DIODE(_05792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13319__A2 (.DIODE(_05807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13335__A1 (.DIODE(_00745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13335__A2 (.DIODE(_02724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13335__B1 (.DIODE(_02728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13335__B2 (.DIODE(_00914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13336__A (.DIODE(_00914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13336__B (.DIODE(_00745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13336__C (.DIODE(_02724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13336__D (.DIODE(_02728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13348__A1 (.DIODE(_01584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13348__A2 (.DIODE(_02306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13348__B1 (.DIODE(_02305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13348__B2 (.DIODE(_01586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13349__A (.DIODE(_01600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13349__B (.DIODE(_01585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13349__C (.DIODE(_02306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13349__D (.DIODE(_02857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13363__A (.DIODE(_00416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13363__B (.DIODE(_01288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13363__C (.DIODE(_02720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13364__A1 (.DIODE(_01289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13364__A2 (.DIODE(_02759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13364__B1 (.DIODE(_02721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13364__B2 (.DIODE(_02008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13365__A1 (.DIODE(_02765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13368__B1 (.DIODE(_02765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13368__B2 (.DIODE(_02008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13376__A1 (.DIODE(_00607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13377__A1 (.DIODE(_01504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13377__B2 (.DIODE(_01508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13378__A (.DIODE(_01664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13378__B (.DIODE(_01505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13389__A2 (.DIODE(_02673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13390__A1 (.DIODE(_00779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13390__A2 (.DIODE(_03681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13390__B1 (.DIODE(_02673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13390__B2 (.DIODE(_01518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13391__A (.DIODE(_01518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13391__B (.DIODE(_01517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13391__C (.DIODE(_03681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13391__D (.DIODE(_02673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13404__A1 (.DIODE(_03414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13404__A2 (.DIODE(_01956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13404__B1 (.DIODE(_03687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13404__B2 (.DIODE(_04714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13405__A (.DIODE(_01066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13405__B (.DIODE(_03414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13405__C (.DIODE(_01955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13405__D (.DIODE(_03686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13410__B1 (.DIODE(_01956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13410__B2 (.DIODE(_04714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13419__A1 (.DIODE(_01183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13419__A2 (.DIODE(_01415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13419__B1 (.DIODE(_01252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13419__B2 (.DIODE(_01108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13420__A (.DIODE(_01061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13420__B (.DIODE(_01181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13420__C (.DIODE(_01414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13420__D (.DIODE(_01250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13430__A_N (.DIODE(_05424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13436__A1 (.DIODE(_05833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13438__A (.DIODE(_03785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13439__A (.DIODE(_01181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13439__B (.DIODE(_01250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13439__C (.DIODE(_02721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13439__D (.DIODE(_02726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13441__A1 (.DIODE(_01250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13441__A2 (.DIODE(_02721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13441__B1 (.DIODE(_02735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13441__B2 (.DIODE(_01182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13442__B (.DIODE(_02765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13443__A2 (.DIODE(_02766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13445__A (.DIODE(_01183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13445__B (.DIODE(_01252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13445__C (.DIODE(_02766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13445__D (.DIODE(_02722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13447__A (.DIODE(_01182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13447__B (.DIODE(_01252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13447__C (.DIODE(_02735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13447__D (.DIODE(_02731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13448__A1 (.DIODE(_01252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13448__A2 (.DIODE(_02736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13448__B1 (.DIODE(_02731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13448__B2 (.DIODE(_01182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13450__B (.DIODE(_02722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13453__A (.DIODE(_03783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13454__B (.DIODE(_02766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13461__A2 (.DIODE(_02722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13462__B (.DIODE(_02735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13463__A1 (.DIODE(_01252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13463__A2 (.DIODE(_02737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13464__A (.DIODE(_01252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13464__C (.DIODE(_02735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13464__D (.DIODE(_02731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13466__B (.DIODE(_02722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13475__A (.DIODE(_02856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13476__A (.DIODE(_01414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13476__C (.DIODE(_01956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13476__D (.DIODE(_03687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13477__A2 (.DIODE(_01956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13477__B1 (.DIODE(_03687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13477__B2 (.DIODE(_01414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13478__C (.DIODE(_01062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13480__A1_N (.DIODE(_01108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13481__A (.DIODE(_01062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13481__B (.DIODE(_01415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13481__C (.DIODE(_01958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13481__D (.DIODE(_03690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13483__A (.DIODE(_02858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13484__C (.DIODE(_01957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13484__D (.DIODE(_03690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13485__A2 (.DIODE(_01957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13485__B1 (.DIODE(_03690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13487__A (.DIODE(_01415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13489__B1 (.DIODE(_01062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13490__A1 (.DIODE(_01062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13496__A1 (.DIODE(_01415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13498__A2 (.DIODE(_03690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13499__C (.DIODE(_03687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13500__C (.DIODE(_01415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13500__D (.DIODE(_03680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13501__A1_N (.DIODE(_01415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13501__A2_N (.DIODE(_03680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13511__A2 (.DIODE(_02722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13512__A2 (.DIODE(_02736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13512__B1 (.DIODE(_02737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13513__C (.DIODE(_02736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13513__D (.DIODE(_02737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13534__A (.DIODE(_02766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13535__A (.DIODE(_01958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13536__A (.DIODE(_02722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13537__A (.DIODE(_03690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13545__B (.DIODE(_02737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13561__B1 (.DIODE(_02736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13561__B2 (.DIODE(_01958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13562__D (.DIODE(_02736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13576__A (.DIODE(_02855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13576__B (.DIODE(_03785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13577__A (.DIODE(_01249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13577__B (.DIODE(_02855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13577__C (.DIODE(_03785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13577__D (.DIODE(_02857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13578__A1 (.DIODE(_01250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13578__A2 (.DIODE(_02858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13580__A (.DIODE(_01414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13580__B (.DIODE(_03783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13582__B (.DIODE(_03785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13582__C (.DIODE(_02858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13582__D (.DIODE(_03783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13583__A1 (.DIODE(_03785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13583__A2 (.DIODE(_02858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13583__B1 (.DIODE(_03783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13583__B2 (.DIODE(_02856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13588__A1 (.DIODE(_01414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13588__A2 (.DIODE(_03783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13590__A (.DIODE(_01181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13590__B (.DIODE(_01250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13590__C (.DIODE(_02856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13590__D (.DIODE(_02858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13591__A1 (.DIODE(_01250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13591__A2 (.DIODE(_02856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13591__B1 (.DIODE(_02858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13591__B2 (.DIODE(_01181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13592__C (.DIODE(_01414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13592__D (.DIODE(_03785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13597__A1 (.DIODE(_01413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13597__A2 (.DIODE(_01249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13597__B1 (.DIODE(_02856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13597__B2 (.DIODE(_01180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13598__A (.DIODE(_01181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13598__B (.DIODE(_01413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13598__C (.DIODE(_01250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13599__A1 (.DIODE(_01061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13599__A2 (.DIODE(_03785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13599__B2 (.DIODE(_02856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13600__A (.DIODE(_01061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13600__B (.DIODE(_03783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13601__A1_N (.DIODE(_01414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13601__A2_N (.DIODE(_03785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13602__A1 (.DIODE(_01061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13602__A2 (.DIODE(_03783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13606__A1 (.DIODE(_02856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13607__A (.DIODE(_01061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13607__B (.DIODE(_03785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13656__A1 (.DIODE(_01252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13656__A2 (.DIODE(_02766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13656__B2 (.DIODE(_01183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13660__A1 (.DIODE(_01415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13660__A2 (.DIODE(_01958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13660__B2 (.DIODE(_01108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13667__A (.DIODE(_01108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13670__A (.DIODE(_01183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13671__A1 (.DIODE(_01183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13671__A2 (.DIODE(_02766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13686__A (.DIODE(_02427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13686__B (.DIODE(_02426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13686__C (.DIODE(_02735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13686__D (.DIODE(_02731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13687__A (.DIODE(_01288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13687__B (.DIODE(_02090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13687__C (.DIODE(_02725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13687__D (.DIODE(_02728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13688__A (.DIODE(_02090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13688__B (.DIODE(_02725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13689__A1 (.DIODE(_01289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13689__A2 (.DIODE(_02730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13691__A (.DIODE(_02088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13691__B (.DIODE(_02720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13692__A1 (.DIODE(_02426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13692__A2 (.DIODE(_02736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13692__B1 (.DIODE(_02737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13692__B2 (.DIODE(_02427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13695__A (.DIODE(_02426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13695__B (.DIODE(_02737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13697__A (.DIODE(_00416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13697__B (.DIODE(_01288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13697__C (.DIODE(_02725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13697__D (.DIODE(_02730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13698__A1 (.DIODE(_01289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13698__A2 (.DIODE(_02726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13698__B1 (.DIODE(_02730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13698__B2 (.DIODE(_01188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13699__C (.DIODE(_02427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13699__D (.DIODE(_02720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13701__A1 (.DIODE(_02426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13701__A2 (.DIODE(_02721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13706__A1 (.DIODE(_01288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13706__A2 (.DIODE(_02720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13706__B1 (.DIODE(_02725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13706__B2 (.DIODE(_00416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13707__A1 (.DIODE(_02726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13708__A (.DIODE(_02427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13708__B (.DIODE(_02759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13710__A (.DIODE(_02759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13711__A1_N (.DIODE(_02427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13711__A2_N (.DIODE(_02721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13713__A1 (.DIODE(_02427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13713__A2 (.DIODE(_02758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13713__B2 (.DIODE(_02726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13714__A (.DIODE(_02426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13714__B (.DIODE(_02759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13715__A1 (.DIODE(_02426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13715__A2 (.DIODE(_02759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13734__A (.DIODE(_00915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13734__B (.DIODE(_02725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13735__A (.DIODE(_00916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13735__B (.DIODE(_02730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13741__A (.DIODE(_02090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13741__B (.DIODE(_02855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13742__A (.DIODE(_02088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13742__B (.DIODE(_02858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13772__A1 (.DIODE(_02765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13798__A (.DIODE(_02188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13798__B (.DIODE(_02190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13798__D (.DIODE(_03680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13799__A (.DIODE(_02187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13799__B (.DIODE(_02189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13799__C (.DIODE(_03686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13799__D (.DIODE(_03683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13800__A (.DIODE(_02187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13800__B (.DIODE(_03682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13801__A1 (.DIODE(_02189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13801__A2 (.DIODE(_03686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13803__A (.DIODE(_03414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13803__B (.DIODE(_03679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13804__A1 (.DIODE(_02190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13804__B1 (.DIODE(_03680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13804__B2 (.DIODE(_02188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13807__A (.DIODE(_02190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13809__A (.DIODE(_02187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13809__B (.DIODE(_02189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13809__C (.DIODE(_01954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13809__D (.DIODE(_03686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13810__A1 (.DIODE(_02189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13810__A2 (.DIODE(_01955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13810__B1 (.DIODE(_03686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13810__B2 (.DIODE(_02188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13811__C (.DIODE(_01400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13811__D (.DIODE(_03683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13813__A1 (.DIODE(_03414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13813__A2 (.DIODE(_03679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13818__A (.DIODE(_01400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13818__B (.DIODE(_02187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13818__C (.DIODE(_03686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13819__A1 (.DIODE(_02187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13819__A2 (.DIODE(_01955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13819__B1 (.DIODE(_03686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13819__B2 (.DIODE(_01400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13820__A1 (.DIODE(_01955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13821__A (.DIODE(_04714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13821__B (.DIODE(_03683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13824__A1_N (.DIODE(_03414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13824__A2_N (.DIODE(_03683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13826__A1 (.DIODE(_00460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13826__A2 (.DIODE(_03683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13826__B2 (.DIODE(_01955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13827__A (.DIODE(_01066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13827__B (.DIODE(_03679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13828__A1 (.DIODE(_04714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13828__A2 (.DIODE(_03680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13847__A (.DIODE(_02189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13847__B (.DIODE(_03783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13853__A (.DIODE(_01517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13853__B (.DIODE(_03679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13958__B (.DIODE(_06540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13969__B (.DIODE(_06552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13970__B (.DIODE(_06540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13981__B (.DIODE(_06552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14022__A (.DIODE(_05424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14025__A1 (.DIODE(_05810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14060__C (.DIODE(_02743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14060__D (.DIODE(_02742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14069__A2 (.DIODE(_02743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14069__B1 (.DIODE(_02742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14070__C (.DIODE(_02743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14070__D (.DIODE(_02742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14074__A4 (.DIODE(_02743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14097__A (.DIODE(_06684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14103__A (.DIODE(_06684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14106__A (.DIODE(_02743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14107__A2 (.DIODE(_02742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14108__B (.DIODE(_02743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14108__D (.DIODE(_02742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14134__A2 (.DIODE(_02742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14134__B2 (.DIODE(_02743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14135__A (.DIODE(_02743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14135__C (.DIODE(_02742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14156__A2 (.DIODE(_05833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14163__A (.DIODE(_02742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14180__A (.DIODE(_02743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14180__C (.DIODE(_02742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14184__A3 (.DIODE(_06778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14196__B (.DIODE(_06778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14201__A (.DIODE(_00344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14201__B (.DIODE(_00410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14211__A (.DIODE(_06800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14212__A1 (.DIODE(_00464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14212__A2 (.DIODE(_02138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14212__B1 (.DIODE(_00344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14212__B2 (.DIODE(_02051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14218__A (.DIODE(_00464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14218__B (.DIODE(_00344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14219__A (.DIODE(_06804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14229__A (.DIODE(_06810_));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap130_A (.DIODE(_05595_));
 sky130_fd_sc_hd__diode_2 ANTENNA_output101_A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_output102_A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_output103_A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_output104_A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_output105_A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_output108_A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_output109_A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_output110_A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_output111_A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_output112_A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_output113_A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_output115_A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_output116_A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_output117_A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_output118_A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_output119_A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_output120_A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_output121_A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_output122_A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_output125_A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_output126_A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_output127_A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_output66_A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_output67_A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_output69_A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_output70_A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_output71_A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_output72_A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_output73_A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_output74_A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_output75_A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_output76_A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_output77_A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_output79_A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_output80_A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_output81_A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_output82_A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_output83_A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_output84_A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_output86_A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_output89_A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_output90_A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_output91_A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_output92_A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_output93_A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_output94_A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_output95_A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_output96_A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_output97_A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_output98_A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_split3_A (.DIODE(_00869_));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_555 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_693 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_704 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_308 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_648 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_678 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_823 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_847 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_366 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_650 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_702 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_680 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_776 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_672 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_644 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_704 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_636 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_791 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_588 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_620 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_702 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_609 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_700 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_711 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_527 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_14 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_560 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_756 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_611 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_703 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_747 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_667 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_650 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_662 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_695 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_535 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_703 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_450 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_415 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_876 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_338 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_508 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_588 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_706 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_676 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_735 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_637 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_664 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_688 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_664 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_676 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_748 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_830 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_859 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_506 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_779 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_860 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_634 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_854 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_507 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_620 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_723 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_675 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_704 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_667 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_722 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_854 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_535 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_855 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_679 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_723 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_777 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_860 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_644 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_702 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_822 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_676 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_728 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_796 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_704 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_802 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_828 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_543 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_859 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_874 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_799 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_622 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_862 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_786 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_790 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_590 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_616 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_646 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_578 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_618 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_786 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_594 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_667 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_702 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_758 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_739 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_779 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_616 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_620 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_646 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_763 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_87 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_871 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_675 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_674 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_832 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_843 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_647 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_683 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_858 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_631 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_588 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_676 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_637 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_591 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_700 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_723 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_762 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_823 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_827 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_395 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_830 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_728 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_738 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_506 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_619 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_650 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_506 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_616 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_846 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_594 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_744 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_812 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_860 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_690 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_718 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_731 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_675 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_594 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_748 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_680 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_788 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_792 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_739 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_693 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_721 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_735 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__clkbuf_4 _07085_ (.A(net33),
    .X(_00300_));
 sky130_fd_sc_hd__buf_4 _07086_ (.A(_00300_),
    .X(_00311_));
 sky130_fd_sc_hd__buf_4 _07087_ (.A(_00311_),
    .X(_00322_));
 sky130_fd_sc_hd__buf_4 _07088_ (.A(_00322_),
    .X(_00333_));
 sky130_fd_sc_hd__buf_6 _07089_ (.A(_00333_),
    .X(_00344_));
 sky130_fd_sc_hd__clkbuf_4 _07090_ (.A(net31),
    .X(_00355_));
 sky130_fd_sc_hd__buf_4 _07091_ (.A(_00355_),
    .X(_00366_));
 sky130_fd_sc_hd__clkbuf_4 _07092_ (.A(_00366_),
    .X(_00377_));
 sky130_fd_sc_hd__buf_4 _07093_ (.A(_00377_),
    .X(_00388_));
 sky130_fd_sc_hd__buf_4 _07094_ (.A(_00388_),
    .X(_00399_));
 sky130_fd_sc_hd__clkbuf_8 _07095_ (.A(_00399_),
    .X(_00410_));
 sky130_fd_sc_hd__buf_6 _07096_ (.A(net1),
    .X(_00420_));
 sky130_fd_sc_hd__clkbuf_4 _07097_ (.A(_00420_),
    .X(_00431_));
 sky130_fd_sc_hd__buf_6 _07098_ (.A(_00431_),
    .X(_00442_));
 sky130_fd_sc_hd__buf_4 _07099_ (.A(_00442_),
    .X(_00453_));
 sky130_fd_sc_hd__buf_4 _07100_ (.A(_00453_),
    .X(_00464_));
 sky130_fd_sc_hd__clkbuf_4 _07101_ (.A(net63),
    .X(_00475_));
 sky130_fd_sc_hd__clkbuf_4 _07102_ (.A(_00475_),
    .X(_00486_));
 sky130_fd_sc_hd__clkbuf_4 _07103_ (.A(_00486_),
    .X(_00497_));
 sky130_fd_sc_hd__buf_4 _07104_ (.A(_00497_),
    .X(_00508_));
 sky130_fd_sc_hd__buf_4 _07105_ (.A(_00508_),
    .X(_00519_));
 sky130_fd_sc_hd__buf_4 _07106_ (.A(_00519_),
    .X(_00530_));
 sky130_fd_sc_hd__clkbuf_4 _07107_ (.A(net29),
    .X(_00541_));
 sky130_fd_sc_hd__nand2_1 _07108_ (.A(_00541_),
    .B(_00300_),
    .Y(_00552_));
 sky130_fd_sc_hd__buf_6 _07109_ (.A(net27),
    .X(_00563_));
 sky130_fd_sc_hd__buf_6 _07110_ (.A(net55),
    .X(_00573_));
 sky130_fd_sc_hd__and4_1 _07111_ (.A(_00563_),
    .B(net28),
    .C(_00573_),
    .D(net44),
    .X(_00584_));
 sky130_fd_sc_hd__a22o_1 _07112_ (.A1(_00563_),
    .A2(_00573_),
    .B1(net44),
    .B2(net28),
    .X(_00595_));
 sky130_fd_sc_hd__and2b_1 _07113_ (.A_N(_00584_),
    .B(_00595_),
    .X(_00606_));
 sky130_fd_sc_hd__xnor2_1 _07114_ (.A(_00552_),
    .B(_00606_),
    .Y(_00617_));
 sky130_fd_sc_hd__clkbuf_4 _07115_ (.A(_00563_),
    .X(_00628_));
 sky130_fd_sc_hd__buf_8 _07116_ (.A(net28),
    .X(_00639_));
 sky130_fd_sc_hd__clkbuf_4 _07117_ (.A(_00639_),
    .X(_00650_));
 sky130_fd_sc_hd__buf_6 _07118_ (.A(net44),
    .X(_00661_));
 sky130_fd_sc_hd__buf_4 _07119_ (.A(_00661_),
    .X(_00672_));
 sky130_fd_sc_hd__and4_1 _07120_ (.A(_00628_),
    .B(_00650_),
    .C(_00672_),
    .D(_00300_),
    .X(_00683_));
 sky130_fd_sc_hd__nand2_1 _07121_ (.A(_00617_),
    .B(_00683_),
    .Y(_00694_));
 sky130_fd_sc_hd__buf_8 _07122_ (.A(net58),
    .X(_00705_));
 sky130_fd_sc_hd__buf_6 _07123_ (.A(net55),
    .X(_00716_));
 sky130_fd_sc_hd__and4_1 _07124_ (.A(net27),
    .B(_00705_),
    .C(net28),
    .D(net161),
    .X(_00726_));
 sky130_fd_sc_hd__a22o_1 _07125_ (.A1(net27),
    .A2(_00705_),
    .B1(net28),
    .B2(_00573_),
    .X(_00737_));
 sky130_fd_sc_hd__and2b_1 _07126_ (.A_N(_00737_),
    .B(_00726_),
    .X(_00748_));
 sky130_fd_sc_hd__nand2_1 _07127_ (.A(_00541_),
    .B(_00661_),
    .Y(_00759_));
 sky130_fd_sc_hd__xnor2_2 _07128_ (.A(_00748_),
    .B(_00759_),
    .Y(_00770_));
 sky130_fd_sc_hd__a31o_1 _07129_ (.A1(net29),
    .A2(net33),
    .A3(_00595_),
    .B1(_00584_),
    .X(_00781_));
 sky130_fd_sc_hd__nand2_1 _07130_ (.A(net30),
    .B(net33),
    .Y(_00792_));
 sky130_fd_sc_hd__xnor2_2 _07131_ (.A(_00781_),
    .B(_00792_),
    .Y(_00803_));
 sky130_fd_sc_hd__xnor2_1 _07132_ (.A(_00770_),
    .B(_00803_),
    .Y(_00814_));
 sky130_fd_sc_hd__nor2_1 _07133_ (.A(_00694_),
    .B(_00814_),
    .Y(_00825_));
 sky130_fd_sc_hd__nand2_1 _07134_ (.A(_00694_),
    .B(_00814_),
    .Y(_00836_));
 sky130_fd_sc_hd__or2b_1 _07135_ (.A(net153),
    .B_N(_00836_),
    .X(_00847_));
 sky130_fd_sc_hd__inv_2 _07136_ (.A(_00847_),
    .Y(_00858_));
 sky130_fd_sc_hd__buf_8 _07137_ (.A(net23),
    .X(_00869_));
 sky130_fd_sc_hd__clkbuf_4 _07138_ (.A(_00869_),
    .X(_00880_));
 sky130_fd_sc_hd__buf_6 _07139_ (.A(_00880_),
    .X(_00891_));
 sky130_fd_sc_hd__clkbuf_4 _07140_ (.A(net59),
    .X(_00901_));
 sky130_fd_sc_hd__nand2_1 _07141_ (.A(_00891_),
    .B(_00901_),
    .Y(_00912_));
 sky130_fd_sc_hd__buf_6 _07142_ (.A(net12),
    .X(_00923_));
 sky130_fd_sc_hd__and4_1 _07143_ (.A(net1),
    .B(_00923_),
    .C(net61),
    .D(net60),
    .X(_00934_));
 sky130_fd_sc_hd__a22o_1 _07144_ (.A1(_00420_),
    .A2(net61),
    .B1(net60),
    .B2(net176),
    .X(_00945_));
 sky130_fd_sc_hd__and2b_1 _07145_ (.A_N(_00934_),
    .B(_00945_),
    .X(_00956_));
 sky130_fd_sc_hd__xnor2_1 _07146_ (.A(_00912_),
    .B(_00956_),
    .Y(_00967_));
 sky130_fd_sc_hd__clkbuf_4 _07147_ (.A(net12),
    .X(_00978_));
 sky130_fd_sc_hd__buf_4 _07148_ (.A(_00978_),
    .X(_00989_));
 sky130_fd_sc_hd__clkbuf_4 _07149_ (.A(net60),
    .X(_01000_));
 sky130_fd_sc_hd__and4_1 _07150_ (.A(_00442_),
    .B(_00989_),
    .C(_01000_),
    .D(_00901_),
    .X(_01011_));
 sky130_fd_sc_hd__nand2_1 _07151_ (.A(_00967_),
    .B(_01011_),
    .Y(_01022_));
 sky130_fd_sc_hd__and4_1 _07152_ (.A(net1),
    .B(net62),
    .C(net12),
    .D(net61),
    .X(_01033_));
 sky130_fd_sc_hd__clkbuf_4 _07153_ (.A(net62),
    .X(_01044_));
 sky130_fd_sc_hd__a22o_1 _07154_ (.A1(net1),
    .A2(_01044_),
    .B1(_00923_),
    .B2(net61),
    .X(_01055_));
 sky130_fd_sc_hd__and2b_1 _07155_ (.A_N(_01033_),
    .B(_01055_),
    .X(_01065_));
 sky130_fd_sc_hd__buf_4 _07156_ (.A(_00869_),
    .X(_01076_));
 sky130_fd_sc_hd__nand2_1 _07157_ (.A(_01076_),
    .B(net60),
    .Y(_01087_));
 sky130_fd_sc_hd__xnor2_2 _07158_ (.A(_01065_),
    .B(_01087_),
    .Y(_01098_));
 sky130_fd_sc_hd__a31o_1 _07159_ (.A1(_00880_),
    .A2(net59),
    .A3(_00945_),
    .B1(_00934_),
    .X(_01109_));
 sky130_fd_sc_hd__clkbuf_4 _07160_ (.A(net26),
    .X(_01120_));
 sky130_fd_sc_hd__nand2_1 _07161_ (.A(_01120_),
    .B(net59),
    .Y(_01131_));
 sky130_fd_sc_hd__xnor2_2 _07162_ (.A(_01109_),
    .B(_01131_),
    .Y(_01142_));
 sky130_fd_sc_hd__xnor2_1 _07163_ (.A(_01098_),
    .B(_01142_),
    .Y(_01153_));
 sky130_fd_sc_hd__nor2_1 _07164_ (.A(_01022_),
    .B(_01153_),
    .Y(_01164_));
 sky130_fd_sc_hd__nand2_1 _07165_ (.A(_01022_),
    .B(_01153_),
    .Y(_01175_));
 sky130_fd_sc_hd__and2b_1 _07166_ (.A_N(net168),
    .B(_01175_),
    .X(_01186_));
 sky130_fd_sc_hd__clkbuf_4 _07167_ (.A(net58),
    .X(_01197_));
 sky130_fd_sc_hd__clkbuf_4 _07168_ (.A(_00716_),
    .X(_01208_));
 sky130_fd_sc_hd__and4_1 _07169_ (.A(_00880_),
    .B(net26),
    .C(_01197_),
    .D(_01208_),
    .X(_01219_));
 sky130_fd_sc_hd__clkbuf_4 _07170_ (.A(net26),
    .X(_01230_));
 sky130_fd_sc_hd__a22o_1 _07171_ (.A1(_00978_),
    .A2(_00705_),
    .B1(_01208_),
    .B2(_00869_),
    .X(_01241_));
 sky130_fd_sc_hd__and4_1 _07172_ (.A(net176),
    .B(net149),
    .C(_00705_),
    .D(_00573_),
    .X(_01251_));
 sky130_fd_sc_hd__a31o_1 _07173_ (.A1(_01230_),
    .A2(_00672_),
    .A3(_01241_),
    .B1(_01251_),
    .X(_01262_));
 sky130_fd_sc_hd__inv_2 _07174_ (.A(_01219_),
    .Y(_01273_));
 sky130_fd_sc_hd__buf_4 _07175_ (.A(_01076_),
    .X(_01284_));
 sky130_fd_sc_hd__clkbuf_4 _07176_ (.A(_01197_),
    .X(_01295_));
 sky130_fd_sc_hd__clkbuf_4 _07177_ (.A(_01208_),
    .X(_01306_));
 sky130_fd_sc_hd__a22o_1 _07178_ (.A1(_01284_),
    .A2(_01295_),
    .B1(_01306_),
    .B2(_01230_),
    .X(_01317_));
 sky130_fd_sc_hd__and3_1 _07179_ (.A(_01262_),
    .B(_01273_),
    .C(_01317_),
    .X(_01328_));
 sky130_fd_sc_hd__clkbuf_4 _07180_ (.A(_01230_),
    .X(_01339_));
 sky130_fd_sc_hd__clkbuf_4 _07181_ (.A(_01339_),
    .X(_01350_));
 sky130_fd_sc_hd__clkbuf_4 _07182_ (.A(_01295_),
    .X(_01361_));
 sky130_fd_sc_hd__buf_4 _07183_ (.A(_00891_),
    .X(_01372_));
 sky130_fd_sc_hd__buf_6 _07184_ (.A(_01372_),
    .X(_01383_));
 sky130_fd_sc_hd__buf_6 _07185_ (.A(_01208_),
    .X(_01394_));
 sky130_fd_sc_hd__buf_4 _07186_ (.A(_01394_),
    .X(_01405_));
 sky130_fd_sc_hd__nand2_1 _07187_ (.A(_01383_),
    .B(_01405_),
    .Y(_01416_));
 sky130_fd_sc_hd__and3_1 _07188_ (.A(_01350_),
    .B(_01361_),
    .C(_01416_),
    .X(_01427_));
 sky130_fd_sc_hd__and2_1 _07189_ (.A(_01328_),
    .B(_01427_),
    .X(_01438_));
 sky130_fd_sc_hd__xor2_2 _07190_ (.A(_01328_),
    .B(_01427_),
    .X(_01448_));
 sky130_fd_sc_hd__or2b_4 _07191_ (.A(_01251_),
    .B_N(_01241_),
    .X(_01459_));
 sky130_fd_sc_hd__buf_4 _07192_ (.A(_00661_),
    .X(_01470_));
 sky130_fd_sc_hd__nand2_1 _07193_ (.A(_01120_),
    .B(_01470_),
    .Y(_01481_));
 sky130_fd_sc_hd__xnor2_2 _07194_ (.A(_01459_),
    .B(_01481_),
    .Y(_01492_));
 sky130_fd_sc_hd__a22o_1 _07195_ (.A1(_00420_),
    .A2(_01197_),
    .B1(_01208_),
    .B2(_00978_),
    .X(_01503_));
 sky130_fd_sc_hd__and4_1 _07196_ (.A(_00420_),
    .B(_00978_),
    .C(_00705_),
    .D(_01208_),
    .X(_01514_));
 sky130_fd_sc_hd__a31o_1 _07197_ (.A1(_01284_),
    .A2(_00672_),
    .A3(_01503_),
    .B1(_01514_),
    .X(_01525_));
 sky130_fd_sc_hd__or2b_4 _07198_ (.A(_01492_),
    .B_N(_01525_),
    .X(_01536_));
 sky130_fd_sc_hd__a21oi_1 _07199_ (.A1(_01273_),
    .A2(_01317_),
    .B1(_01262_),
    .Y(_01547_));
 sky130_fd_sc_hd__nor2_1 _07200_ (.A(_01328_),
    .B(_01547_),
    .Y(_01558_));
 sky130_fd_sc_hd__xor2_2 _07201_ (.A(_01536_),
    .B(_01558_),
    .X(_01569_));
 sky130_fd_sc_hd__nand2_1 _07202_ (.A(_01230_),
    .B(_00300_),
    .Y(_01580_));
 sky130_fd_sc_hd__a22o_1 _07203_ (.A1(_00420_),
    .A2(_01208_),
    .B1(_00661_),
    .B2(_00978_),
    .X(_01591_));
 sky130_fd_sc_hd__and4_1 _07204_ (.A(_00420_),
    .B(_00978_),
    .C(_01208_),
    .D(net44),
    .X(_01602_));
 sky130_fd_sc_hd__a31o_1 _07205_ (.A1(_01076_),
    .A2(net33),
    .A3(_01591_),
    .B1(_01602_),
    .X(_01613_));
 sky130_fd_sc_hd__or2b_1 _07206_ (.A(_01580_),
    .B_N(_01613_),
    .X(_01624_));
 sky130_fd_sc_hd__and2b_1 _07207_ (.A_N(_01514_),
    .B(_01503_),
    .X(_01635_));
 sky130_fd_sc_hd__nand2_1 _07208_ (.A(_00891_),
    .B(_00672_),
    .Y(_01645_));
 sky130_fd_sc_hd__xnor2_1 _07209_ (.A(_01635_),
    .B(_01645_),
    .Y(_01656_));
 sky130_fd_sc_hd__xnor2_2 _07210_ (.A(_01613_),
    .B(_01580_),
    .Y(_01667_));
 sky130_fd_sc_hd__nand2_1 _07211_ (.A(_01656_),
    .B(_01667_),
    .Y(_01678_));
 sky130_fd_sc_hd__xor2_1 _07212_ (.A(_01525_),
    .B(_01492_),
    .X(_01689_));
 sky130_fd_sc_hd__nand3_2 _07213_ (.A(_01624_),
    .B(_01678_),
    .C(_01689_),
    .Y(_01700_));
 sky130_fd_sc_hd__and2b_1 _07214_ (.A_N(_01602_),
    .B(_01591_),
    .X(_01711_));
 sky130_fd_sc_hd__nand2_1 _07215_ (.A(_01284_),
    .B(_00300_),
    .Y(_01722_));
 sky130_fd_sc_hd__xnor2_1 _07216_ (.A(_01711_),
    .B(_01722_),
    .Y(_01733_));
 sky130_fd_sc_hd__buf_4 _07217_ (.A(_00672_),
    .X(_01744_));
 sky130_fd_sc_hd__and4_2 _07218_ (.A(_00442_),
    .B(_00989_),
    .C(_01744_),
    .D(_00311_),
    .X(_01755_));
 sky130_fd_sc_hd__nand2_1 _07219_ (.A(_01733_),
    .B(_01755_),
    .Y(_01766_));
 sky130_fd_sc_hd__xnor2_1 _07220_ (.A(_01656_),
    .B(_01667_),
    .Y(_01777_));
 sky130_fd_sc_hd__nor2_4 _07221_ (.A(_01766_),
    .B(_01777_),
    .Y(_01788_));
 sky130_fd_sc_hd__a21o_1 _07222_ (.A1(_01624_),
    .A2(_01678_),
    .B1(_01689_),
    .X(_01799_));
 sky130_fd_sc_hd__a21boi_4 _07223_ (.A1(_01700_),
    .A2(_01788_),
    .B1_N(_01799_),
    .Y(_01810_));
 sky130_fd_sc_hd__and2b_1 _07224_ (.A_N(_01536_),
    .B(_01558_),
    .X(_01821_));
 sky130_fd_sc_hd__o21bai_4 _07225_ (.A1(_01569_),
    .A2(_01810_),
    .B1_N(_01821_),
    .Y(_01832_));
 sky130_fd_sc_hd__and2_4 _07226_ (.A(_01448_),
    .B(_01832_),
    .X(_01842_));
 sky130_fd_sc_hd__or4_4 _07227_ (.A(_01186_),
    .B(_01219_),
    .C(_01438_),
    .D(_01842_),
    .X(_01853_));
 sky130_fd_sc_hd__o31ai_1 _07228_ (.A1(_01219_),
    .A2(_01438_),
    .A3(_01842_),
    .B1(_01186_),
    .Y(_01864_));
 sky130_fd_sc_hd__nand2_1 _07229_ (.A(_01853_),
    .B(_01864_),
    .Y(_01875_));
 sky130_fd_sc_hd__xnor2_2 _07230_ (.A(_00858_),
    .B(_01875_),
    .Y(_01886_));
 sky130_fd_sc_hd__or2_1 _07231_ (.A(_00967_),
    .B(_01011_),
    .X(_01897_));
 sky130_fd_sc_hd__nand2_1 _07232_ (.A(_01022_),
    .B(_01897_),
    .Y(_01908_));
 sky130_fd_sc_hd__xnor2_2 _07233_ (.A(_01448_),
    .B(_01832_),
    .Y(_01919_));
 sky130_fd_sc_hd__nand2_1 _07234_ (.A(_01908_),
    .B(_01919_),
    .Y(_01930_));
 sky130_fd_sc_hd__or2_1 _07235_ (.A(_00617_),
    .B(_00683_),
    .X(_01941_));
 sky130_fd_sc_hd__nand2_1 _07236_ (.A(_00694_),
    .B(_01941_),
    .Y(_01952_));
 sky130_fd_sc_hd__o21ai_1 _07237_ (.A1(_01908_),
    .A2(_01919_),
    .B1(_01952_),
    .Y(_01963_));
 sky130_fd_sc_hd__nand2_1 _07238_ (.A(_01930_),
    .B(_01963_),
    .Y(_01974_));
 sky130_fd_sc_hd__xnor2_1 _07239_ (.A(_01886_),
    .B(_01974_),
    .Y(_01985_));
 sky130_fd_sc_hd__buf_4 _07240_ (.A(_01000_),
    .X(_01996_));
 sky130_fd_sc_hd__buf_4 _07241_ (.A(_01996_),
    .X(_02007_));
 sky130_fd_sc_hd__clkbuf_4 _07242_ (.A(_02007_),
    .X(_02018_));
 sky130_fd_sc_hd__buf_4 _07243_ (.A(_00901_),
    .X(_02029_));
 sky130_fd_sc_hd__buf_4 _07244_ (.A(_02029_),
    .X(_02040_));
 sky130_fd_sc_hd__buf_4 _07245_ (.A(_00989_),
    .X(_02051_));
 sky130_fd_sc_hd__a22oi_2 _07246_ (.A1(_00442_),
    .A2(_02018_),
    .B1(_02040_),
    .B2(_02051_),
    .Y(_02061_));
 sky130_fd_sc_hd__nor2_1 _07247_ (.A(_01011_),
    .B(_02061_),
    .Y(_02072_));
 sky130_fd_sc_hd__xor2_2 _07248_ (.A(_01569_),
    .B(net181),
    .X(_02083_));
 sky130_fd_sc_hd__nor2_1 _07249_ (.A(_02072_),
    .B(net184),
    .Y(_02094_));
 sky130_fd_sc_hd__clkbuf_4 _07250_ (.A(_00628_),
    .X(_02105_));
 sky130_fd_sc_hd__clkbuf_4 _07251_ (.A(_02105_),
    .X(_02116_));
 sky130_fd_sc_hd__clkbuf_4 _07252_ (.A(_00672_),
    .X(_02127_));
 sky130_fd_sc_hd__buf_4 _07253_ (.A(_02127_),
    .X(_02138_));
 sky130_fd_sc_hd__clkbuf_4 _07254_ (.A(_00650_),
    .X(_02149_));
 sky130_fd_sc_hd__buf_2 _07255_ (.A(_02149_),
    .X(_02160_));
 sky130_fd_sc_hd__buf_4 _07256_ (.A(_02160_),
    .X(_02171_));
 sky130_fd_sc_hd__a22oi_1 _07257_ (.A1(_02116_),
    .A2(_02138_),
    .B1(_00333_),
    .B2(_02171_),
    .Y(_02182_));
 sky130_fd_sc_hd__or2_1 _07258_ (.A(_00683_),
    .B(_02182_),
    .X(_02193_));
 sky130_fd_sc_hd__nand2_1 _07259_ (.A(_02072_),
    .B(net184),
    .Y(_02204_));
 sky130_fd_sc_hd__o21ai_1 _07260_ (.A1(_02094_),
    .A2(_02193_),
    .B1(_02204_),
    .Y(_02215_));
 sky130_fd_sc_hd__xor2_1 _07261_ (.A(_01908_),
    .B(_01919_),
    .X(_02226_));
 sky130_fd_sc_hd__xnor2_1 _07262_ (.A(_01952_),
    .B(_02226_),
    .Y(_02237_));
 sky130_fd_sc_hd__or2_1 _07263_ (.A(_02215_),
    .B(_02237_),
    .X(_02248_));
 sky130_fd_sc_hd__buf_4 _07264_ (.A(_02116_),
    .X(_02259_));
 sky130_fd_sc_hd__and2_2 _07265_ (.A(_02259_),
    .B(_00333_),
    .X(_02270_));
 sky130_fd_sc_hd__clkbuf_4 _07266_ (.A(_02040_),
    .X(_02280_));
 sky130_fd_sc_hd__and3_1 _07267_ (.A(_01799_),
    .B(_01700_),
    .C(_01788_),
    .X(_02291_));
 sky130_fd_sc_hd__a21oi_1 _07268_ (.A1(net156),
    .A2(_01700_),
    .B1(_01788_),
    .Y(_02302_));
 sky130_fd_sc_hd__nor2_1 _07269_ (.A(_02291_),
    .B(_02302_),
    .Y(_02313_));
 sky130_fd_sc_hd__and3_1 _07270_ (.A(_00453_),
    .B(_02280_),
    .C(_02313_),
    .X(_02324_));
 sky130_fd_sc_hd__clkbuf_4 _07271_ (.A(_02280_),
    .X(_02335_));
 sky130_fd_sc_hd__a21o_1 _07272_ (.A1(_00453_),
    .A2(_02335_),
    .B1(_02313_),
    .X(_02346_));
 sky130_fd_sc_hd__o21a_1 _07273_ (.A1(_02270_),
    .A2(_02324_),
    .B1(_02346_),
    .X(_02357_));
 sky130_fd_sc_hd__xnor2_1 _07274_ (.A(_02072_),
    .B(_02083_),
    .Y(_02368_));
 sky130_fd_sc_hd__xnor2_1 _07275_ (.A(_02193_),
    .B(_02368_),
    .Y(_02379_));
 sky130_fd_sc_hd__inv_2 _07276_ (.A(_02379_),
    .Y(_02390_));
 sky130_fd_sc_hd__and2_1 _07277_ (.A(_02357_),
    .B(_02390_),
    .X(_02401_));
 sky130_fd_sc_hd__and2_1 _07278_ (.A(_02215_),
    .B(_02237_),
    .X(_02412_));
 sky130_fd_sc_hd__a21o_2 _07279_ (.A1(_02248_),
    .A2(_02401_),
    .B1(_02412_),
    .X(_02423_));
 sky130_fd_sc_hd__and3_1 _07280_ (.A(_01886_),
    .B(_01930_),
    .C(_01963_),
    .X(_02434_));
 sky130_fd_sc_hd__a21o_1 _07281_ (.A1(_01985_),
    .A2(_02423_),
    .B1(_02434_),
    .X(_02445_));
 sky130_fd_sc_hd__buf_4 _07282_ (.A(_02335_),
    .X(_02456_));
 sky130_fd_sc_hd__clkbuf_8 _07283_ (.A(_02259_),
    .X(_02467_));
 sky130_fd_sc_hd__nand2_1 _07284_ (.A(_02456_),
    .B(_02467_),
    .Y(_02478_));
 sky130_fd_sc_hd__nand2_1 _07285_ (.A(_00847_),
    .B(_01864_),
    .Y(_02489_));
 sky130_fd_sc_hd__or2b_1 _07286_ (.A(_01131_),
    .B_N(_01109_),
    .X(_02499_));
 sky130_fd_sc_hd__nand2_1 _07287_ (.A(_01098_),
    .B(_01142_),
    .Y(_02510_));
 sky130_fd_sc_hd__a31o_1 _07288_ (.A1(_00891_),
    .A2(_01000_),
    .A3(_01055_),
    .B1(_01033_),
    .X(_02521_));
 sky130_fd_sc_hd__and4_1 _07289_ (.A(net62),
    .B(net12),
    .C(net61),
    .D(_00869_),
    .X(_02532_));
 sky130_fd_sc_hd__a22o_1 _07290_ (.A1(net62),
    .A2(_00923_),
    .B1(net61),
    .B2(_00869_),
    .X(_02543_));
 sky130_fd_sc_hd__and2b_1 _07291_ (.A_N(_02532_),
    .B(_02543_),
    .X(_02554_));
 sky130_fd_sc_hd__nand2_1 _07292_ (.A(net60),
    .B(net26),
    .Y(_02565_));
 sky130_fd_sc_hd__xnor2_1 _07293_ (.A(_02554_),
    .B(_02565_),
    .Y(_02576_));
 sky130_fd_sc_hd__xnor2_2 _07294_ (.A(_02521_),
    .B(net152),
    .Y(_02587_));
 sky130_fd_sc_hd__a21oi_2 _07295_ (.A1(_02499_),
    .A2(_02510_),
    .B1(_02587_),
    .Y(_02598_));
 sky130_fd_sc_hd__nand3_1 _07296_ (.A(_02499_),
    .B(_02510_),
    .C(_02587_),
    .Y(_02609_));
 sky130_fd_sc_hd__and2b_1 _07297_ (.A_N(_02598_),
    .B(_02609_),
    .X(_02620_));
 sky130_fd_sc_hd__xnor2_1 _07298_ (.A(net169),
    .B(_02620_),
    .Y(_02631_));
 sky130_fd_sc_hd__or2b_1 _07299_ (.A(_00792_),
    .B_N(_00781_),
    .X(_02642_));
 sky130_fd_sc_hd__nand2_1 _07300_ (.A(_00770_),
    .B(_00803_),
    .Y(_02653_));
 sky130_fd_sc_hd__clkbuf_4 _07301_ (.A(net29),
    .X(_02664_));
 sky130_fd_sc_hd__a31o_1 _07302_ (.A1(_02664_),
    .A2(_00672_),
    .A3(_00737_),
    .B1(_00726_),
    .X(_02675_));
 sky130_fd_sc_hd__and4_1 _07303_ (.A(_00705_),
    .B(net28),
    .C(_00573_),
    .D(net29),
    .X(_02686_));
 sky130_fd_sc_hd__a22o_1 _07304_ (.A1(_00705_),
    .A2(_00639_),
    .B1(_00573_),
    .B2(net29),
    .X(_02697_));
 sky130_fd_sc_hd__and2b_1 _07305_ (.A_N(_02686_),
    .B(_02697_),
    .X(_02708_));
 sky130_fd_sc_hd__clkbuf_4 _07306_ (.A(net30),
    .X(_02719_));
 sky130_fd_sc_hd__nand2_1 _07307_ (.A(_01470_),
    .B(_02719_),
    .Y(_02729_));
 sky130_fd_sc_hd__xnor2_2 _07308_ (.A(_02708_),
    .B(_02729_),
    .Y(_02740_));
 sky130_fd_sc_hd__xnor2_2 _07309_ (.A(_02675_),
    .B(_02740_),
    .Y(_02751_));
 sky130_fd_sc_hd__a21oi_1 _07310_ (.A1(_02642_),
    .A2(_02653_),
    .B1(_02751_),
    .Y(_02762_));
 sky130_fd_sc_hd__nand3_2 _07311_ (.A(_02642_),
    .B(_02653_),
    .C(_02751_),
    .Y(_02773_));
 sky130_fd_sc_hd__and2b_1 _07312_ (.A_N(_02762_),
    .B(_02773_),
    .X(_02784_));
 sky130_fd_sc_hd__xnor2_1 _07313_ (.A(net153),
    .B(_02784_),
    .Y(_02795_));
 sky130_fd_sc_hd__nor2_1 _07314_ (.A(_02631_),
    .B(_02795_),
    .Y(_02806_));
 sky130_fd_sc_hd__and2_1 _07315_ (.A(_02631_),
    .B(_02795_),
    .X(_02817_));
 sky130_fd_sc_hd__nor2_1 _07316_ (.A(_02806_),
    .B(_02817_),
    .Y(_02828_));
 sky130_fd_sc_hd__a21oi_1 _07317_ (.A1(_01853_),
    .A2(_02489_),
    .B1(_02828_),
    .Y(_02839_));
 sky130_fd_sc_hd__o31a_1 _07318_ (.A1(_01219_),
    .A2(_01438_),
    .A3(_01842_),
    .B1(_01186_),
    .X(_02850_));
 sky130_fd_sc_hd__o211a_1 _07319_ (.A1(_00858_),
    .A2(_02850_),
    .B1(_02828_),
    .C1(_01853_),
    .X(_02861_));
 sky130_fd_sc_hd__nor2_1 _07320_ (.A(_02839_),
    .B(_02861_),
    .Y(_02872_));
 sky130_fd_sc_hd__xnor2_2 _07321_ (.A(_02478_),
    .B(_02872_),
    .Y(_02883_));
 sky130_fd_sc_hd__nand2_2 _07322_ (.A(_02445_),
    .B(_02883_),
    .Y(_02894_));
 sky130_fd_sc_hd__or2_1 _07323_ (.A(_02445_),
    .B(_02883_),
    .X(_02905_));
 sky130_fd_sc_hd__and2_1 _07324_ (.A(_02894_),
    .B(_02905_),
    .X(_02916_));
 sky130_fd_sc_hd__a21o_1 _07325_ (.A1(_00464_),
    .A2(_00530_),
    .B1(_02916_),
    .X(_02927_));
 sky130_fd_sc_hd__and3_1 _07326_ (.A(_00464_),
    .B(_00530_),
    .C(_02916_),
    .X(_02938_));
 sky130_fd_sc_hd__a31o_1 _07327_ (.A1(_00344_),
    .A2(_00410_),
    .A3(_02927_),
    .B1(_02938_),
    .X(_02949_));
 sky130_fd_sc_hd__buf_4 _07328_ (.A(net32),
    .X(_02960_));
 sky130_fd_sc_hd__clkbuf_4 _07329_ (.A(_02960_),
    .X(_02971_));
 sky130_fd_sc_hd__buf_4 _07330_ (.A(_02971_),
    .X(_02982_));
 sky130_fd_sc_hd__clkbuf_4 _07331_ (.A(_02982_),
    .X(_02993_));
 sky130_fd_sc_hd__clkbuf_4 _07332_ (.A(_02993_),
    .X(_03004_));
 sky130_fd_sc_hd__buf_4 _07333_ (.A(_03004_),
    .X(_03015_));
 sky130_fd_sc_hd__a22oi_2 _07334_ (.A1(_02138_),
    .A2(_00410_),
    .B1(_03015_),
    .B2(_00333_),
    .Y(_03026_));
 sky130_fd_sc_hd__and4_1 _07335_ (.A(_01470_),
    .B(net33),
    .C(_00355_),
    .D(_02971_),
    .X(_03037_));
 sky130_fd_sc_hd__nor2_1 _07336_ (.A(_03026_),
    .B(_03037_),
    .Y(_03048_));
 sky130_fd_sc_hd__clkbuf_4 _07337_ (.A(_02018_),
    .X(_03059_));
 sky130_fd_sc_hd__clkbuf_4 _07338_ (.A(_03059_),
    .X(_03070_));
 sky130_fd_sc_hd__a22o_1 _07339_ (.A1(_03070_),
    .A2(_02259_),
    .B1(_02171_),
    .B2(_02280_),
    .X(_03081_));
 sky130_fd_sc_hd__and4_1 _07340_ (.A(_02007_),
    .B(_02029_),
    .C(_02105_),
    .D(_02149_),
    .X(_03092_));
 sky130_fd_sc_hd__inv_2 _07341_ (.A(_03092_),
    .Y(_03103_));
 sky130_fd_sc_hd__and2_1 _07342_ (.A(_03081_),
    .B(_03103_),
    .X(_03114_));
 sky130_fd_sc_hd__nand2_1 _07343_ (.A(_02576_),
    .B(_02521_),
    .Y(_03125_));
 sky130_fd_sc_hd__a31o_1 _07344_ (.A1(net60),
    .A2(net26),
    .A3(_02543_),
    .B1(_02532_),
    .X(_03136_));
 sky130_fd_sc_hd__buf_2 _07345_ (.A(net61),
    .X(_03147_));
 sky130_fd_sc_hd__a22o_1 _07346_ (.A1(_01044_),
    .A2(_00880_),
    .B1(net26),
    .B2(_03147_),
    .X(_03158_));
 sky130_fd_sc_hd__nand4_1 _07347_ (.A(_01044_),
    .B(_03147_),
    .C(_00880_),
    .D(net26),
    .Y(_03169_));
 sky130_fd_sc_hd__nand2_1 _07348_ (.A(_03158_),
    .B(_03169_),
    .Y(_03180_));
 sky130_fd_sc_hd__xor2_1 _07349_ (.A(_03136_),
    .B(_03180_),
    .X(_03191_));
 sky130_fd_sc_hd__nor2_1 _07350_ (.A(_03125_),
    .B(_03191_),
    .Y(_03202_));
 sky130_fd_sc_hd__and2_4 _07351_ (.A(_03125_),
    .B(_03191_),
    .X(_03213_));
 sky130_fd_sc_hd__or2_4 _07352_ (.A(_03202_),
    .B(_03213_),
    .X(_03224_));
 sky130_fd_sc_hd__a21oi_2 _07353_ (.A1(_01164_),
    .A2(_02609_),
    .B1(_02598_),
    .Y(_03235_));
 sky130_fd_sc_hd__xor2_2 _07354_ (.A(_03224_),
    .B(net147),
    .X(_03246_));
 sky130_fd_sc_hd__nand2_1 _07355_ (.A(_02675_),
    .B(net189),
    .Y(_03257_));
 sky130_fd_sc_hd__buf_4 _07356_ (.A(_02719_),
    .X(_03268_));
 sky130_fd_sc_hd__a31o_1 _07357_ (.A1(_01744_),
    .A2(_03268_),
    .A3(_02697_),
    .B1(_02686_),
    .X(_03279_));
 sky130_fd_sc_hd__a22o_1 _07358_ (.A1(_01295_),
    .A2(_02664_),
    .B1(_02719_),
    .B2(_01306_),
    .X(_03290_));
 sky130_fd_sc_hd__nand4_2 _07359_ (.A(_01295_),
    .B(_01405_),
    .C(_02664_),
    .D(_02719_),
    .Y(_03301_));
 sky130_fd_sc_hd__nand2_1 _07360_ (.A(_03290_),
    .B(_03301_),
    .Y(_03312_));
 sky130_fd_sc_hd__xor2_1 _07361_ (.A(_03279_),
    .B(_03312_),
    .X(_03323_));
 sky130_fd_sc_hd__nor2_1 _07362_ (.A(_03257_),
    .B(_03323_),
    .Y(_03334_));
 sky130_fd_sc_hd__nand2_1 _07363_ (.A(_03257_),
    .B(_03323_),
    .Y(_03345_));
 sky130_fd_sc_hd__or2b_1 _07364_ (.A(_03334_),
    .B_N(_03345_),
    .X(_03356_));
 sky130_fd_sc_hd__a21o_1 _07365_ (.A1(_00825_),
    .A2(_02773_),
    .B1(_02762_),
    .X(_03367_));
 sky130_fd_sc_hd__xnor2_2 _07366_ (.A(_03356_),
    .B(net188),
    .Y(_03378_));
 sky130_fd_sc_hd__xor2_1 _07367_ (.A(_03246_),
    .B(_03378_),
    .X(_03389_));
 sky130_fd_sc_hd__and2_4 _07368_ (.A(_02806_),
    .B(_03389_),
    .X(_03400_));
 sky130_fd_sc_hd__or2_4 _07369_ (.A(_02806_),
    .B(_03389_),
    .X(_03411_));
 sky130_fd_sc_hd__and2b_1 _07370_ (.A_N(_03400_),
    .B(_03411_),
    .X(_03422_));
 sky130_fd_sc_hd__xnor2_2 _07371_ (.A(_03114_),
    .B(_03422_),
    .Y(_03433_));
 sky130_fd_sc_hd__a21oi_2 _07372_ (.A1(_02456_),
    .A2(_02467_),
    .B1(_02861_),
    .Y(_03444_));
 sky130_fd_sc_hd__nor3_2 _07373_ (.A(_02839_),
    .B(_03433_),
    .C(_03444_),
    .Y(_03455_));
 sky130_fd_sc_hd__o21a_1 _07374_ (.A1(_02839_),
    .A2(_03444_),
    .B1(_03433_),
    .X(_03466_));
 sky130_fd_sc_hd__nor2_4 _07375_ (.A(_03466_),
    .B(_03455_),
    .Y(_03477_));
 sky130_fd_sc_hd__xor2_4 _07376_ (.A(_02894_),
    .B(_03477_),
    .X(_03488_));
 sky130_fd_sc_hd__clkbuf_4 _07377_ (.A(net64),
    .X(_03499_));
 sky130_fd_sc_hd__clkbuf_4 _07378_ (.A(_03499_),
    .X(_03510_));
 sky130_fd_sc_hd__clkbuf_4 _07379_ (.A(_03510_),
    .X(_03521_));
 sky130_fd_sc_hd__clkbuf_4 _07380_ (.A(_03521_),
    .X(_03532_));
 sky130_fd_sc_hd__clkbuf_4 _07381_ (.A(_03532_),
    .X(_03543_));
 sky130_fd_sc_hd__buf_4 _07382_ (.A(_03543_),
    .X(_03554_));
 sky130_fd_sc_hd__a22oi_2 _07383_ (.A1(_00453_),
    .A2(_03554_),
    .B1(_00519_),
    .B2(_02051_),
    .Y(_03565_));
 sky130_fd_sc_hd__buf_4 _07384_ (.A(_00431_),
    .X(_03576_));
 sky130_fd_sc_hd__clkbuf_4 _07385_ (.A(_00978_),
    .X(_03587_));
 sky130_fd_sc_hd__and4_1 _07386_ (.A(_03576_),
    .B(_03587_),
    .C(_03499_),
    .D(net63),
    .X(_03598_));
 sky130_fd_sc_hd__or2_2 _07387_ (.A(_03565_),
    .B(_03598_),
    .X(_03609_));
 sky130_fd_sc_hd__xnor2_1 _07388_ (.A(_03488_),
    .B(_03609_),
    .Y(_03620_));
 sky130_fd_sc_hd__xnor2_2 _07389_ (.A(_03048_),
    .B(_03620_),
    .Y(_03631_));
 sky130_fd_sc_hd__nand2_2 _07390_ (.A(_02949_),
    .B(_03631_),
    .Y(_03642_));
 sky130_fd_sc_hd__or2_1 _07391_ (.A(_02949_),
    .B(_03631_),
    .X(_03653_));
 sky130_fd_sc_hd__and2_1 _07392_ (.A(_03642_),
    .B(_03653_),
    .X(_03664_));
 sky130_fd_sc_hd__clkbuf_1 _07393_ (.A(_03664_),
    .X(net128));
 sky130_fd_sc_hd__buf_6 _07394_ (.A(net8),
    .X(_03685_));
 sky130_fd_sc_hd__clkbuf_4 _07395_ (.A(_03685_),
    .X(_03696_));
 sky130_fd_sc_hd__buf_4 _07396_ (.A(_03696_),
    .X(_03707_));
 sky130_fd_sc_hd__buf_4 _07397_ (.A(net9),
    .X(_03718_));
 sky130_fd_sc_hd__clkbuf_4 _07398_ (.A(_03718_),
    .X(_03729_));
 sky130_fd_sc_hd__buf_4 _07399_ (.A(_03729_),
    .X(_03740_));
 sky130_fd_sc_hd__and4_1 _07400_ (.A(_02127_),
    .B(_00322_),
    .C(_03707_),
    .D(_03740_),
    .X(_03751_));
 sky130_fd_sc_hd__clkbuf_4 _07401_ (.A(net10),
    .X(_03762_));
 sky130_fd_sc_hd__clkbuf_4 _07402_ (.A(_03762_),
    .X(_03773_));
 sky130_fd_sc_hd__nand2_1 _07403_ (.A(_00322_),
    .B(_03773_),
    .Y(_03784_));
 sky130_fd_sc_hd__and4_1 _07404_ (.A(_01394_),
    .B(_01470_),
    .C(_03685_),
    .D(_03718_),
    .X(_03795_));
 sky130_fd_sc_hd__a22o_1 _07405_ (.A1(_01394_),
    .A2(_03685_),
    .B1(_03718_),
    .B2(_01470_),
    .X(_03806_));
 sky130_fd_sc_hd__and2b_1 _07406_ (.A_N(_03795_),
    .B(_03806_),
    .X(_03817_));
 sky130_fd_sc_hd__xnor2_1 _07407_ (.A(_03784_),
    .B(_03817_),
    .Y(_03828_));
 sky130_fd_sc_hd__nand2_1 _07408_ (.A(_03751_),
    .B(_03828_),
    .Y(_03839_));
 sky130_fd_sc_hd__buf_2 _07409_ (.A(_01197_),
    .X(_03850_));
 sky130_fd_sc_hd__and4_1 _07410_ (.A(_03850_),
    .B(_01394_),
    .C(net8),
    .D(_03718_),
    .X(_03861_));
 sky130_fd_sc_hd__a22o_1 _07411_ (.A1(_03850_),
    .A2(_03685_),
    .B1(_03718_),
    .B2(_01306_),
    .X(_03872_));
 sky130_fd_sc_hd__and2b_1 _07412_ (.A_N(_03861_),
    .B(_03872_),
    .X(_03883_));
 sky130_fd_sc_hd__clkbuf_4 _07413_ (.A(net10),
    .X(_03894_));
 sky130_fd_sc_hd__nand2_1 _07414_ (.A(_02127_),
    .B(_03894_),
    .Y(_03905_));
 sky130_fd_sc_hd__xnor2_1 _07415_ (.A(_03883_),
    .B(_03905_),
    .Y(_03916_));
 sky130_fd_sc_hd__a31o_1 _07416_ (.A1(_00311_),
    .A2(_03762_),
    .A3(_03806_),
    .B1(_03795_),
    .X(_03927_));
 sky130_fd_sc_hd__clkbuf_4 _07417_ (.A(net11),
    .X(_03938_));
 sky130_fd_sc_hd__nand2_1 _07418_ (.A(_00311_),
    .B(_03938_),
    .Y(_03949_));
 sky130_fd_sc_hd__xnor2_1 _07419_ (.A(_03927_),
    .B(_03949_),
    .Y(_03960_));
 sky130_fd_sc_hd__xnor2_1 _07420_ (.A(_03916_),
    .B(_03960_),
    .Y(_03971_));
 sky130_fd_sc_hd__nor2_1 _07421_ (.A(_03839_),
    .B(_03971_),
    .Y(_03982_));
 sky130_fd_sc_hd__nand2_1 _07422_ (.A(_03839_),
    .B(_03971_),
    .Y(_03993_));
 sky130_fd_sc_hd__or2b_4 _07423_ (.A(_03982_),
    .B_N(_03993_),
    .X(_04004_));
 sky130_fd_sc_hd__buf_2 _07424_ (.A(net41),
    .X(_04015_));
 sky130_fd_sc_hd__clkbuf_4 _07425_ (.A(_04015_),
    .X(_04026_));
 sky130_fd_sc_hd__clkbuf_4 _07426_ (.A(_04026_),
    .X(_04037_));
 sky130_fd_sc_hd__clkbuf_4 _07427_ (.A(net40),
    .X(_04048_));
 sky130_fd_sc_hd__clkbuf_4 _07428_ (.A(_04048_),
    .X(_04059_));
 sky130_fd_sc_hd__and4_1 _07429_ (.A(_00442_),
    .B(_02051_),
    .C(_04037_),
    .D(_04059_),
    .X(_04070_));
 sky130_fd_sc_hd__clkbuf_4 _07430_ (.A(_01284_),
    .X(_04081_));
 sky130_fd_sc_hd__nand2_1 _07431_ (.A(_04081_),
    .B(_04048_),
    .Y(_04092_));
 sky130_fd_sc_hd__clkbuf_4 _07432_ (.A(net42),
    .X(_04103_));
 sky130_fd_sc_hd__and4_1 _07433_ (.A(_03576_),
    .B(_03587_),
    .C(_04015_),
    .D(_04103_),
    .X(_04114_));
 sky130_fd_sc_hd__a22o_1 _07434_ (.A1(_03587_),
    .A2(_04015_),
    .B1(_04103_),
    .B2(_03576_),
    .X(_04125_));
 sky130_fd_sc_hd__and2b_1 _07435_ (.A_N(_04114_),
    .B(_04125_),
    .X(_04136_));
 sky130_fd_sc_hd__xnor2_1 _07436_ (.A(_04092_),
    .B(_04136_),
    .Y(_04147_));
 sky130_fd_sc_hd__nand2_1 _07437_ (.A(_04070_),
    .B(_04147_),
    .Y(_04158_));
 sky130_fd_sc_hd__buf_2 _07438_ (.A(_00978_),
    .X(_04169_));
 sky130_fd_sc_hd__buf_2 _07439_ (.A(net42),
    .X(_04180_));
 sky130_fd_sc_hd__buf_4 _07440_ (.A(net43),
    .X(_04191_));
 sky130_fd_sc_hd__and4_1 _07441_ (.A(_00431_),
    .B(_04169_),
    .C(_04180_),
    .D(_04191_),
    .X(_04202_));
 sky130_fd_sc_hd__a22o_1 _07442_ (.A1(_03587_),
    .A2(_04103_),
    .B1(_04191_),
    .B2(_03576_),
    .X(_04213_));
 sky130_fd_sc_hd__and2b_1 _07443_ (.A_N(_04202_),
    .B(_04213_),
    .X(_04224_));
 sky130_fd_sc_hd__nand2_1 _07444_ (.A(_01372_),
    .B(_04026_),
    .Y(_04235_));
 sky130_fd_sc_hd__xnor2_1 _07445_ (.A(_04224_),
    .B(_04235_),
    .Y(_04246_));
 sky130_fd_sc_hd__a31o_1 _07446_ (.A1(_01284_),
    .A2(net40),
    .A3(_04125_),
    .B1(_04114_),
    .X(_04257_));
 sky130_fd_sc_hd__clkbuf_4 _07447_ (.A(_01230_),
    .X(_04268_));
 sky130_fd_sc_hd__nand2_1 _07448_ (.A(_04268_),
    .B(_04048_),
    .Y(_04279_));
 sky130_fd_sc_hd__xnor2_1 _07449_ (.A(_04257_),
    .B(_04279_),
    .Y(_04290_));
 sky130_fd_sc_hd__xnor2_1 _07450_ (.A(_04246_),
    .B(_04290_),
    .Y(_04301_));
 sky130_fd_sc_hd__nor2_1 _07451_ (.A(_04158_),
    .B(_04301_),
    .Y(_04312_));
 sky130_fd_sc_hd__nand2_1 _07452_ (.A(_04158_),
    .B(_04301_),
    .Y(_04323_));
 sky130_fd_sc_hd__nand2b_2 _07453_ (.A_N(_04312_),
    .B(_04323_),
    .Y(_04334_));
 sky130_fd_sc_hd__nand4_2 _07454_ (.A(_01996_),
    .B(_00901_),
    .C(_00366_),
    .D(_02982_),
    .Y(_04345_));
 sky130_fd_sc_hd__a22o_1 _07455_ (.A1(_02018_),
    .A2(_00388_),
    .B1(_03004_),
    .B2(_02040_),
    .X(_04356_));
 sky130_fd_sc_hd__buf_6 _07456_ (.A(net2),
    .X(_04367_));
 sky130_fd_sc_hd__buf_4 _07457_ (.A(_04367_),
    .X(_04378_));
 sky130_fd_sc_hd__a22o_1 _07458_ (.A1(net58),
    .A2(net31),
    .B1(net32),
    .B2(net175),
    .X(_04389_));
 sky130_fd_sc_hd__and4_1 _07459_ (.A(net58),
    .B(net163),
    .C(net31),
    .D(net32),
    .X(_04400_));
 sky130_fd_sc_hd__a31o_1 _07460_ (.A1(_01470_),
    .A2(_04378_),
    .A3(_04389_),
    .B1(net164),
    .X(_04411_));
 sky130_fd_sc_hd__and4_1 _07461_ (.A(net58),
    .B(net175),
    .C(net32),
    .D(net2),
    .X(_04422_));
 sky130_fd_sc_hd__a22o_1 _07462_ (.A1(net58),
    .A2(net32),
    .B1(net2),
    .B2(net163),
    .X(_04433_));
 sky130_fd_sc_hd__and2b_1 _07463_ (.A_N(_04422_),
    .B(_04433_),
    .X(_04444_));
 sky130_fd_sc_hd__buf_2 _07464_ (.A(net3),
    .X(_04455_));
 sky130_fd_sc_hd__nand2_1 _07465_ (.A(_00661_),
    .B(_04455_),
    .Y(_04466_));
 sky130_fd_sc_hd__xnor2_1 _07466_ (.A(_04444_),
    .B(_04466_),
    .Y(_04477_));
 sky130_fd_sc_hd__a31o_1 _07467_ (.A1(_00661_),
    .A2(_04455_),
    .A3(_04433_),
    .B1(_04422_),
    .X(_04488_));
 sky130_fd_sc_hd__nand4_2 _07468_ (.A(_03850_),
    .B(_01394_),
    .C(_04378_),
    .D(_04455_),
    .Y(_04499_));
 sky130_fd_sc_hd__buf_2 _07469_ (.A(_00573_),
    .X(_04510_));
 sky130_fd_sc_hd__a22o_1 _07470_ (.A1(_01197_),
    .A2(_04367_),
    .B1(_04455_),
    .B2(_04510_),
    .X(_04521_));
 sky130_fd_sc_hd__and3_2 _07471_ (.A(_04488_),
    .B(_04499_),
    .C(_04521_),
    .X(_04532_));
 sky130_fd_sc_hd__a21oi_1 _07472_ (.A1(_04499_),
    .A2(_04521_),
    .B1(_04488_),
    .Y(_04543_));
 sky130_fd_sc_hd__nor2_1 _07473_ (.A(_04532_),
    .B(_04543_),
    .Y(_04554_));
 sky130_fd_sc_hd__and3_1 _07474_ (.A(_04411_),
    .B(_04477_),
    .C(_04554_),
    .X(_04565_));
 sky130_fd_sc_hd__a21oi_1 _07475_ (.A1(_04411_),
    .A2(_04477_),
    .B1(_04554_),
    .Y(_04576_));
 sky130_fd_sc_hd__nor2_1 _07476_ (.A(_04565_),
    .B(_04576_),
    .Y(_04587_));
 sky130_fd_sc_hd__buf_4 _07477_ (.A(_04455_),
    .X(_04598_));
 sky130_fd_sc_hd__a22o_1 _07478_ (.A1(net163),
    .A2(net31),
    .B1(net32),
    .B2(net44),
    .X(_04609_));
 sky130_fd_sc_hd__and4_1 _07479_ (.A(net162),
    .B(net44),
    .C(net31),
    .D(net32),
    .X(_04620_));
 sky130_fd_sc_hd__a31o_1 _07480_ (.A1(net33),
    .A2(_04367_),
    .A3(_04609_),
    .B1(_04620_),
    .X(_04631_));
 sky130_fd_sc_hd__and3_1 _07481_ (.A(_00300_),
    .B(_04598_),
    .C(_04631_),
    .X(_04642_));
 sky130_fd_sc_hd__or2b_1 _07482_ (.A(_04400_),
    .B_N(_04389_),
    .X(_04653_));
 sky130_fd_sc_hd__nand2_1 _07483_ (.A(_00661_),
    .B(_04367_),
    .Y(_04664_));
 sky130_fd_sc_hd__xnor2_1 _07484_ (.A(_04653_),
    .B(_04664_),
    .Y(_04675_));
 sky130_fd_sc_hd__nand2_1 _07485_ (.A(net33),
    .B(_04455_),
    .Y(_04686_));
 sky130_fd_sc_hd__xnor2_1 _07486_ (.A(_04631_),
    .B(_04686_),
    .Y(_04697_));
 sky130_fd_sc_hd__and2b_1 _07487_ (.A_N(_04697_),
    .B(_04675_),
    .X(_04708_));
 sky130_fd_sc_hd__xor2_1 _07488_ (.A(_04411_),
    .B(_04477_),
    .X(_04719_));
 sky130_fd_sc_hd__or3_4 _07489_ (.A(_04642_),
    .B(_04708_),
    .C(_04719_),
    .X(_04730_));
 sky130_fd_sc_hd__nand2_1 _07490_ (.A(net33),
    .B(_04367_),
    .Y(_04741_));
 sky130_fd_sc_hd__and2b_1 _07491_ (.A_N(_04620_),
    .B(_04609_),
    .X(_04752_));
 sky130_fd_sc_hd__xnor2_1 _07492_ (.A(_04741_),
    .B(_04752_),
    .Y(_04763_));
 sky130_fd_sc_hd__and2_1 _07493_ (.A(_03037_),
    .B(_04763_),
    .X(_04774_));
 sky130_fd_sc_hd__xnor2_1 _07494_ (.A(net154),
    .B(net170),
    .Y(_04785_));
 sky130_fd_sc_hd__and2_2 _07495_ (.A(_04774_),
    .B(_04785_),
    .X(_04796_));
 sky130_fd_sc_hd__o21a_1 _07496_ (.A1(_04642_),
    .A2(_04708_),
    .B1(_04719_),
    .X(_04807_));
 sky130_fd_sc_hd__a21oi_1 _07497_ (.A1(_04730_),
    .A2(_04796_),
    .B1(_04807_),
    .Y(_04818_));
 sky130_fd_sc_hd__xnor2_1 _07498_ (.A(_04587_),
    .B(_04818_),
    .Y(_04829_));
 sky130_fd_sc_hd__a21oi_1 _07499_ (.A1(_04345_),
    .A2(_04356_),
    .B1(_04829_),
    .Y(_04840_));
 sky130_fd_sc_hd__clkbuf_4 _07500_ (.A(net5),
    .X(_04851_));
 sky130_fd_sc_hd__clkbuf_4 _07501_ (.A(_04851_),
    .X(_04862_));
 sky130_fd_sc_hd__buf_4 _07502_ (.A(net4),
    .X(_04873_));
 sky130_fd_sc_hd__nand4_2 _07503_ (.A(_01744_),
    .B(_00311_),
    .C(_04862_),
    .D(_04873_),
    .Y(_04884_));
 sky130_fd_sc_hd__clkbuf_4 _07504_ (.A(_04862_),
    .X(_04895_));
 sky130_fd_sc_hd__clkbuf_4 _07505_ (.A(_04895_),
    .X(_04906_));
 sky130_fd_sc_hd__clkbuf_4 _07506_ (.A(_04906_),
    .X(_04917_));
 sky130_fd_sc_hd__clkbuf_4 _07507_ (.A(_04873_),
    .X(_04928_));
 sky130_fd_sc_hd__buf_4 _07508_ (.A(_04928_),
    .X(_04939_));
 sky130_fd_sc_hd__a22o_1 _07509_ (.A1(_00333_),
    .A2(_04917_),
    .B1(_04939_),
    .B2(_02138_),
    .X(_04950_));
 sky130_fd_sc_hd__nand2_2 _07510_ (.A(_04884_),
    .B(_04950_),
    .Y(_04961_));
 sky130_fd_sc_hd__and3_1 _07511_ (.A(_04345_),
    .B(_04356_),
    .C(_04829_),
    .X(_04972_));
 sky130_fd_sc_hd__o21bai_2 _07512_ (.A1(_04840_),
    .A2(_04961_),
    .B1_N(_04972_),
    .Y(_04983_));
 sky130_fd_sc_hd__and4_1 _07513_ (.A(_00573_),
    .B(net44),
    .C(_04851_),
    .D(net4),
    .X(_04994_));
 sky130_fd_sc_hd__a22o_1 _07514_ (.A1(net44),
    .A2(_04851_),
    .B1(net4),
    .B2(_00573_),
    .X(_05005_));
 sky130_fd_sc_hd__or2b_1 _07515_ (.A(_04994_),
    .B_N(_05005_),
    .X(_05016_));
 sky130_fd_sc_hd__clkbuf_4 _07516_ (.A(net6),
    .X(_05027_));
 sky130_fd_sc_hd__nand2_1 _07517_ (.A(_00300_),
    .B(_05027_),
    .Y(_05038_));
 sky130_fd_sc_hd__xnor2_1 _07518_ (.A(_05016_),
    .B(_05038_),
    .Y(_05049_));
 sky130_fd_sc_hd__or2_1 _07519_ (.A(_04884_),
    .B(_05049_),
    .X(_05060_));
 sky130_fd_sc_hd__nand2_1 _07520_ (.A(_04884_),
    .B(_05049_),
    .Y(_05071_));
 sky130_fd_sc_hd__and2_1 _07521_ (.A(_05060_),
    .B(_05071_),
    .X(_05082_));
 sky130_fd_sc_hd__and4_1 _07522_ (.A(_03147_),
    .B(net60),
    .C(_00355_),
    .D(_02960_),
    .X(_05093_));
 sky130_fd_sc_hd__a22o_1 _07523_ (.A1(_03147_),
    .A2(_00355_),
    .B1(_02960_),
    .B2(net60),
    .X(_05104_));
 sky130_fd_sc_hd__and4b_1 _07524_ (.A_N(_05093_),
    .B(_05104_),
    .C(_00901_),
    .D(_04378_),
    .X(_05115_));
 sky130_fd_sc_hd__inv_2 _07525_ (.A(_05104_),
    .Y(_05126_));
 sky130_fd_sc_hd__o2bb2a_1 _07526_ (.A1_N(_00901_),
    .A2_N(_04378_),
    .B1(_05093_),
    .B2(_05126_),
    .X(_05137_));
 sky130_fd_sc_hd__or3_4 _07527_ (.A(_04345_),
    .B(_05115_),
    .C(_05137_),
    .X(_05148_));
 sky130_fd_sc_hd__o21ai_1 _07528_ (.A1(_05115_),
    .A2(_05137_),
    .B1(_04345_),
    .Y(_05159_));
 sky130_fd_sc_hd__nand2_1 _07529_ (.A(_05148_),
    .B(_05159_),
    .Y(_05170_));
 sky130_fd_sc_hd__buf_4 _07530_ (.A(_04598_),
    .X(_05181_));
 sky130_fd_sc_hd__clkbuf_4 _07531_ (.A(_04378_),
    .X(_05192_));
 sky130_fd_sc_hd__buf_4 _07532_ (.A(_05192_),
    .X(_05203_));
 sky130_fd_sc_hd__nand2_1 _07533_ (.A(_01405_),
    .B(_05203_),
    .Y(_05214_));
 sky130_fd_sc_hd__and3_1 _07534_ (.A(_01361_),
    .B(_05181_),
    .C(_05214_),
    .X(_05225_));
 sky130_fd_sc_hd__xnor2_2 _07535_ (.A(_04532_),
    .B(_05225_),
    .Y(_05236_));
 sky130_fd_sc_hd__a21o_1 _07536_ (.A1(_04730_),
    .A2(_04796_),
    .B1(_04807_),
    .X(_05247_));
 sky130_fd_sc_hd__a21o_1 _07537_ (.A1(_04587_),
    .A2(_05247_),
    .B1(_04565_),
    .X(_05258_));
 sky130_fd_sc_hd__xor2_2 _07538_ (.A(_05236_),
    .B(_05258_),
    .X(_05269_));
 sky130_fd_sc_hd__xnor2_1 _07539_ (.A(_05170_),
    .B(_05269_),
    .Y(_05280_));
 sky130_fd_sc_hd__xnor2_2 _07540_ (.A(_05082_),
    .B(_05280_),
    .Y(_05291_));
 sky130_fd_sc_hd__xnor2_1 _07541_ (.A(_04983_),
    .B(_05291_),
    .Y(_05302_));
 sky130_fd_sc_hd__and2_2 _07542_ (.A(_00333_),
    .B(_04939_),
    .X(_05313_));
 sky130_fd_sc_hd__or2b_1 _07543_ (.A(_04807_),
    .B_N(_04730_),
    .X(_05324_));
 sky130_fd_sc_hd__xnor2_2 _07544_ (.A(_05324_),
    .B(_04796_),
    .Y(_05335_));
 sky130_fd_sc_hd__and3_1 _07545_ (.A(_02335_),
    .B(_00399_),
    .C(_05335_),
    .X(_05346_));
 sky130_fd_sc_hd__a21o_1 _07546_ (.A1(_02456_),
    .A2(_00399_),
    .B1(_05335_),
    .X(_05357_));
 sky130_fd_sc_hd__o21ai_2 _07547_ (.A1(_05313_),
    .A2(_05346_),
    .B1(_05357_),
    .Y(_05368_));
 sky130_fd_sc_hd__or2_1 _07548_ (.A(_04972_),
    .B(_04840_),
    .X(_05379_));
 sky130_fd_sc_hd__xnor2_2 _07549_ (.A(_04961_),
    .B(_05379_),
    .Y(_05390_));
 sky130_fd_sc_hd__nor2_1 _07550_ (.A(_05368_),
    .B(_05390_),
    .Y(_05401_));
 sky130_fd_sc_hd__xnor2_1 _07551_ (.A(_05302_),
    .B(_05401_),
    .Y(_05412_));
 sky130_fd_sc_hd__o21ba_4 _07552_ (.A1(_03224_),
    .A2(_03235_),
    .B1_N(_03202_),
    .X(_05423_));
 sky130_fd_sc_hd__and3_1 _07553_ (.A(_03136_),
    .B(_03158_),
    .C(_03169_),
    .X(_05434_));
 sky130_fd_sc_hd__clkbuf_4 _07554_ (.A(_01044_),
    .X(_05445_));
 sky130_fd_sc_hd__buf_4 _07555_ (.A(_05445_),
    .X(_05456_));
 sky130_fd_sc_hd__clkbuf_4 _07556_ (.A(_03147_),
    .X(_05467_));
 sky130_fd_sc_hd__buf_4 _07557_ (.A(_05467_),
    .X(_05478_));
 sky130_fd_sc_hd__nand2_1 _07558_ (.A(_05478_),
    .B(_01383_),
    .Y(_05489_));
 sky130_fd_sc_hd__and3_1 _07559_ (.A(_05456_),
    .B(_01350_),
    .C(_05489_),
    .X(_05500_));
 sky130_fd_sc_hd__xor2_2 _07560_ (.A(_05434_),
    .B(_05500_),
    .X(_05511_));
 sky130_fd_sc_hd__and2b_1 _07561_ (.A_N(_05511_),
    .B(_05423_),
    .X(_05522_));
 sky130_fd_sc_hd__a21bo_1 _07562_ (.A1(_05434_),
    .A2(_05500_),
    .B1_N(_03169_),
    .X(_05533_));
 sky130_fd_sc_hd__a21oi_2 _07563_ (.A1(_03345_),
    .A2(_03367_),
    .B1(_03334_),
    .Y(_05544_));
 sky130_fd_sc_hd__and3_1 _07564_ (.A(_03279_),
    .B(_03290_),
    .C(_03301_),
    .X(_05555_));
 sky130_fd_sc_hd__buf_4 _07565_ (.A(_03268_),
    .X(_05566_));
 sky130_fd_sc_hd__clkbuf_4 _07566_ (.A(_02664_),
    .X(_05577_));
 sky130_fd_sc_hd__buf_4 _07567_ (.A(_05577_),
    .X(_05588_));
 sky130_fd_sc_hd__nand2_1 _07568_ (.A(_01405_),
    .B(_05588_),
    .Y(_05599_));
 sky130_fd_sc_hd__and3_1 _07569_ (.A(_01361_),
    .B(_05566_),
    .C(_05599_),
    .X(_05610_));
 sky130_fd_sc_hd__xor2_2 _07570_ (.A(_05555_),
    .B(_05610_),
    .X(_05621_));
 sky130_fd_sc_hd__and2b_1 _07571_ (.A_N(_05621_),
    .B(_05544_),
    .X(_05632_));
 sky130_fd_sc_hd__a21bo_1 _07572_ (.A1(_05555_),
    .A2(_05610_),
    .B1_N(_03301_),
    .X(_05643_));
 sky130_fd_sc_hd__o22ai_4 _07573_ (.A1(net151),
    .A2(_05533_),
    .B1(_05632_),
    .B2(_05643_),
    .Y(_05654_));
 sky130_fd_sc_hd__or4_4 _07574_ (.A(_05522_),
    .B(_05533_),
    .C(_05632_),
    .D(_05643_),
    .X(_05665_));
 sky130_fd_sc_hd__xnor2_2 _07575_ (.A(_05621_),
    .B(_05544_),
    .Y(_05676_));
 sky130_fd_sc_hd__xnor2_2 _07576_ (.A(_05511_),
    .B(net190),
    .Y(_05687_));
 sky130_fd_sc_hd__and2_1 _07577_ (.A(_05676_),
    .B(_05687_),
    .X(_05698_));
 sky130_fd_sc_hd__a21oi_2 _07578_ (.A1(_05654_),
    .A2(_05665_),
    .B1(_05698_),
    .Y(_05709_));
 sky130_fd_sc_hd__and3_1 _07579_ (.A(_05654_),
    .B(_05698_),
    .C(_05665_),
    .X(_05720_));
 sky130_fd_sc_hd__clkbuf_4 _07580_ (.A(_03147_),
    .X(_05731_));
 sky130_fd_sc_hd__clkbuf_4 _07581_ (.A(_00639_),
    .X(_05742_));
 sky130_fd_sc_hd__and4_1 _07582_ (.A(_05731_),
    .B(_01000_),
    .C(_00628_),
    .D(_05742_),
    .X(_05753_));
 sky130_fd_sc_hd__a22o_1 _07583_ (.A1(_05731_),
    .A2(_00628_),
    .B1(_05742_),
    .B2(_01000_),
    .X(_05761_));
 sky130_fd_sc_hd__and4b_1 _07584_ (.A_N(_05753_),
    .B(_05761_),
    .C(_00901_),
    .D(_02664_),
    .X(_05771_));
 sky130_fd_sc_hd__inv_2 _07585_ (.A(_05761_),
    .Y(_05780_));
 sky130_fd_sc_hd__o2bb2a_1 _07586_ (.A1_N(_02029_),
    .A2_N(_05588_),
    .B1(_05753_),
    .B2(_05780_),
    .X(_05790_));
 sky130_fd_sc_hd__or2_1 _07587_ (.A(_05771_),
    .B(_05790_),
    .X(_05800_));
 sky130_fd_sc_hd__or2_1 _07588_ (.A(_03103_),
    .B(_05800_),
    .X(_05808_));
 sky130_fd_sc_hd__and4_1 _07589_ (.A(_05445_),
    .B(_05467_),
    .C(_02105_),
    .D(_00650_),
    .X(_05818_));
 sky130_fd_sc_hd__a22o_1 _07590_ (.A1(_05456_),
    .A2(_02105_),
    .B1(_00650_),
    .B2(_05467_),
    .X(_05827_));
 sky130_fd_sc_hd__and2b_1 _07591_ (.A_N(_05818_),
    .B(_05827_),
    .X(_05837_));
 sky130_fd_sc_hd__nand2_1 _07592_ (.A(_02007_),
    .B(_05588_),
    .Y(_05847_));
 sky130_fd_sc_hd__xnor2_1 _07593_ (.A(_05837_),
    .B(_05847_),
    .Y(_05857_));
 sky130_fd_sc_hd__o211ai_2 _07594_ (.A1(_05753_),
    .A2(_05771_),
    .B1(_02029_),
    .C1(_05566_),
    .Y(_05868_));
 sky130_fd_sc_hd__a211o_1 _07595_ (.A1(_02029_),
    .A2(_05566_),
    .B1(_05753_),
    .C1(_05771_),
    .X(_05879_));
 sky130_fd_sc_hd__and2_1 _07596_ (.A(_05868_),
    .B(_05879_),
    .X(_05890_));
 sky130_fd_sc_hd__nand2_1 _07597_ (.A(_05857_),
    .B(_05890_),
    .Y(_05901_));
 sky130_fd_sc_hd__or2_1 _07598_ (.A(_05857_),
    .B(_05890_),
    .X(_05912_));
 sky130_fd_sc_hd__nand2_1 _07599_ (.A(_05901_),
    .B(_05912_),
    .Y(_05923_));
 sky130_fd_sc_hd__nor2_1 _07600_ (.A(_05808_),
    .B(_05923_),
    .Y(_05934_));
 sky130_fd_sc_hd__and2_1 _07601_ (.A(_05808_),
    .B(_05923_),
    .X(_05945_));
 sky130_fd_sc_hd__nor2_1 _07602_ (.A(_05934_),
    .B(_05945_),
    .Y(_05956_));
 sky130_fd_sc_hd__o21ai_2 _07603_ (.A1(_05709_),
    .A2(_05720_),
    .B1(_05956_),
    .Y(_05967_));
 sky130_fd_sc_hd__a31o_1 _07604_ (.A1(_05654_),
    .A2(_05698_),
    .A3(_05665_),
    .B1(_05956_),
    .X(_05977_));
 sky130_fd_sc_hd__or2_4 _07605_ (.A(_05709_),
    .B(_05977_),
    .X(_05988_));
 sky130_fd_sc_hd__nand2_2 _07606_ (.A(net191),
    .B(net192),
    .Y(_05999_));
 sky130_fd_sc_hd__xnor2_2 _07607_ (.A(_05676_),
    .B(_05687_),
    .Y(_06010_));
 sky130_fd_sc_hd__nand2_1 _07608_ (.A(_03103_),
    .B(_05800_),
    .Y(_06021_));
 sky130_fd_sc_hd__nand2_2 _07609_ (.A(_05808_),
    .B(_06021_),
    .Y(_06032_));
 sky130_fd_sc_hd__o21a_1 _07610_ (.A1(_05999_),
    .A2(_06010_),
    .B1(_06032_),
    .X(_06043_));
 sky130_fd_sc_hd__a21o_1 _07611_ (.A1(_05999_),
    .A2(_06010_),
    .B1(_06043_),
    .X(_06054_));
 sky130_fd_sc_hd__a21oi_2 _07612_ (.A1(_05967_),
    .A2(_05988_),
    .B1(_06054_),
    .Y(_06065_));
 sky130_fd_sc_hd__nand3_4 _07613_ (.A(net187),
    .B(_05988_),
    .C(_06054_),
    .Y(_06076_));
 sky130_fd_sc_hd__xor2_2 _07614_ (.A(_05999_),
    .B(_06010_),
    .X(_06087_));
 sky130_fd_sc_hd__xnor2_4 _07615_ (.A(_06032_),
    .B(_06087_),
    .Y(_06098_));
 sky130_fd_sc_hd__a21o_1 _07616_ (.A1(_03114_),
    .A2(_03411_),
    .B1(_03400_),
    .X(_06109_));
 sky130_fd_sc_hd__xor2_4 _07617_ (.A(_06098_),
    .B(_06109_),
    .X(_06120_));
 sky130_fd_sc_hd__nand3b_4 _07618_ (.A_N(_06065_),
    .B(_06076_),
    .C(_06120_),
    .Y(_06131_));
 sky130_fd_sc_hd__nand4b_4 _07619_ (.A_N(_06131_),
    .B(_02883_),
    .C(_02445_),
    .D(_03477_),
    .Y(_06142_));
 sky130_fd_sc_hd__and2_1 _07620_ (.A(_06098_),
    .B(_06109_),
    .X(_06153_));
 sky130_fd_sc_hd__a21o_1 _07621_ (.A1(net140),
    .A2(_06120_),
    .B1(_06153_),
    .X(_06164_));
 sky130_fd_sc_hd__a21oi_4 _07622_ (.A1(_06076_),
    .A2(_06164_),
    .B1(net183),
    .Y(_06175_));
 sky130_fd_sc_hd__a31o_1 _07623_ (.A1(_02007_),
    .A2(_05588_),
    .A3(_05827_),
    .B1(_05818_),
    .X(_06186_));
 sky130_fd_sc_hd__and4_1 _07624_ (.A(_05445_),
    .B(_05467_),
    .C(_05742_),
    .D(_02664_),
    .X(_06197_));
 sky130_fd_sc_hd__nand2_1 _07625_ (.A(_05467_),
    .B(_00541_),
    .Y(_06208_));
 sky130_fd_sc_hd__a21boi_1 _07626_ (.A1(_05445_),
    .A2(_00650_),
    .B1_N(_06208_),
    .Y(_06219_));
 sky130_fd_sc_hd__and4bb_1 _07627_ (.A_N(_06197_),
    .B_N(_06219_),
    .C(_01996_),
    .D(_03268_),
    .X(_06230_));
 sky130_fd_sc_hd__o2bb2a_1 _07628_ (.A1_N(_02007_),
    .A2_N(_05566_),
    .B1(_06197_),
    .B2(_06219_),
    .X(_06241_));
 sky130_fd_sc_hd__nor2_1 _07629_ (.A(_06230_),
    .B(_06241_),
    .Y(_06252_));
 sky130_fd_sc_hd__and2_1 _07630_ (.A(_06186_),
    .B(_06252_),
    .X(_06263_));
 sky130_fd_sc_hd__nor2_1 _07631_ (.A(_06186_),
    .B(_06252_),
    .Y(_06274_));
 sky130_fd_sc_hd__or2_1 _07632_ (.A(_06263_),
    .B(_06274_),
    .X(_06285_));
 sky130_fd_sc_hd__a21oi_1 _07633_ (.A1(_05868_),
    .A2(_05901_),
    .B1(_06285_),
    .Y(_06296_));
 sky130_fd_sc_hd__and3_1 _07634_ (.A(_05868_),
    .B(_05901_),
    .C(_06285_),
    .X(_06307_));
 sky130_fd_sc_hd__nor2_1 _07635_ (.A(_06296_),
    .B(_06307_),
    .Y(_06318_));
 sky130_fd_sc_hd__xnor2_1 _07636_ (.A(_05934_),
    .B(_06318_),
    .Y(_06329_));
 sky130_fd_sc_hd__nor2_1 _07637_ (.A(_05654_),
    .B(_06329_),
    .Y(_06340_));
 sky130_fd_sc_hd__and2_1 _07638_ (.A(_05654_),
    .B(_06329_),
    .X(_06351_));
 sky130_fd_sc_hd__or2_1 _07639_ (.A(_06340_),
    .B(_06351_),
    .X(_06362_));
 sky130_fd_sc_hd__or2b_1 _07640_ (.A(_05709_),
    .B_N(_05977_),
    .X(_06373_));
 sky130_fd_sc_hd__nor2_1 _07641_ (.A(_06362_),
    .B(_06373_),
    .Y(_06384_));
 sky130_fd_sc_hd__nand2_1 _07642_ (.A(_06362_),
    .B(_06373_),
    .Y(_06395_));
 sky130_fd_sc_hd__or2b_1 _07643_ (.A(_06384_),
    .B_N(_06395_),
    .X(_06406_));
 sky130_fd_sc_hd__clkbuf_4 _07644_ (.A(_05456_),
    .X(_06417_));
 sky130_fd_sc_hd__buf_4 _07645_ (.A(_06417_),
    .X(_06428_));
 sky130_fd_sc_hd__clkbuf_4 _07646_ (.A(_05478_),
    .X(_06439_));
 sky130_fd_sc_hd__clkbuf_4 _07647_ (.A(_06439_),
    .X(_06450_));
 sky130_fd_sc_hd__clkbuf_4 _07648_ (.A(_05588_),
    .X(_06461_));
 sky130_fd_sc_hd__clkbuf_4 _07649_ (.A(_06461_),
    .X(_06472_));
 sky130_fd_sc_hd__clkbuf_4 _07650_ (.A(_05566_),
    .X(_06483_));
 sky130_fd_sc_hd__buf_4 _07651_ (.A(_06483_),
    .X(_06494_));
 sky130_fd_sc_hd__nand4_2 _07652_ (.A(_06428_),
    .B(_06450_),
    .C(_06472_),
    .D(_06494_),
    .Y(_06505_));
 sky130_fd_sc_hd__a22o_1 _07653_ (.A1(_06428_),
    .A2(_06472_),
    .B1(_06483_),
    .B2(_06439_),
    .X(_06516_));
 sky130_fd_sc_hd__o211a_2 _07654_ (.A1(_06197_),
    .A2(_06230_),
    .B1(_06505_),
    .C1(_06516_),
    .X(_06527_));
 sky130_fd_sc_hd__a211oi_1 _07655_ (.A1(_06505_),
    .A2(_06516_),
    .B1(_06197_),
    .C1(_06230_),
    .Y(_06538_));
 sky130_fd_sc_hd__nor2_1 _07656_ (.A(_06527_),
    .B(_06538_),
    .Y(_06549_));
 sky130_fd_sc_hd__xnor2_1 _07657_ (.A(_06263_),
    .B(_06549_),
    .Y(_06560_));
 sky130_fd_sc_hd__a21oi_1 _07658_ (.A1(_05934_),
    .A2(_06318_),
    .B1(_06296_),
    .Y(_06571_));
 sky130_fd_sc_hd__nor2_1 _07659_ (.A(_06560_),
    .B(_06571_),
    .Y(_06582_));
 sky130_fd_sc_hd__and2_1 _07660_ (.A(_06560_),
    .B(_06571_),
    .X(_06593_));
 sky130_fd_sc_hd__nor2_1 _07661_ (.A(_06582_),
    .B(_06593_),
    .Y(_06604_));
 sky130_fd_sc_hd__xnor2_1 _07662_ (.A(_06604_),
    .B(_06340_),
    .Y(_06615_));
 sky130_fd_sc_hd__clkbuf_4 _07663_ (.A(_06428_),
    .X(_06626_));
 sky130_fd_sc_hd__buf_4 _07664_ (.A(_06494_),
    .X(_06637_));
 sky130_fd_sc_hd__and3_1 _07665_ (.A(_06626_),
    .B(_06637_),
    .C(_06208_),
    .X(_06648_));
 sky130_fd_sc_hd__xor2_2 _07666_ (.A(_06527_),
    .B(_06648_),
    .X(_06658_));
 sky130_fd_sc_hd__a21o_1 _07667_ (.A1(_06263_),
    .A2(_06549_),
    .B1(_06582_),
    .X(_06669_));
 sky130_fd_sc_hd__xnor2_2 _07668_ (.A(_06658_),
    .B(_06669_),
    .Y(_06680_));
 sky130_fd_sc_hd__a2111oi_4 _07669_ (.A1(_06142_),
    .A2(_06175_),
    .B1(_06406_),
    .C1(_06615_),
    .D1(_06680_),
    .Y(_06691_));
 sky130_fd_sc_hd__o21ai_1 _07670_ (.A1(_06340_),
    .A2(_06384_),
    .B1(_06604_),
    .Y(_06701_));
 sky130_fd_sc_hd__nor2_1 _07671_ (.A(_06680_),
    .B(_06701_),
    .Y(_06712_));
 sky130_fd_sc_hd__nor2_1 _07672_ (.A(_06712_),
    .B(net179),
    .Y(_06723_));
 sky130_fd_sc_hd__clkbuf_4 _07673_ (.A(net37),
    .X(_06733_));
 sky130_fd_sc_hd__clkbuf_4 _07674_ (.A(net36),
    .X(_06744_));
 sky130_fd_sc_hd__and4_1 _07675_ (.A(_00442_),
    .B(_00989_),
    .C(_06733_),
    .D(_06744_),
    .X(_06755_));
 sky130_fd_sc_hd__buf_4 _07676_ (.A(_06733_),
    .X(_06765_));
 sky130_fd_sc_hd__buf_4 _07677_ (.A(_06744_),
    .X(_06775_));
 sky130_fd_sc_hd__a22oi_1 _07678_ (.A1(_00442_),
    .A2(_06765_),
    .B1(_06775_),
    .B2(_02051_),
    .Y(_06785_));
 sky130_fd_sc_hd__nor2_1 _07679_ (.A(_06755_),
    .B(_06785_),
    .Y(_06790_));
 sky130_fd_sc_hd__a22o_1 _07680_ (.A1(net1),
    .A2(net35),
    .B1(net34),
    .B2(net12),
    .X(_06797_));
 sky130_fd_sc_hd__and4_1 _07681_ (.A(net1),
    .B(net12),
    .C(net35),
    .D(net34),
    .X(_06802_));
 sky130_fd_sc_hd__a31o_1 _07682_ (.A1(_01076_),
    .A2(_03499_),
    .A3(_06797_),
    .B1(_06802_),
    .X(_06809_));
 sky130_fd_sc_hd__and4_1 _07683_ (.A(net12),
    .B(net23),
    .C(net35),
    .D(net34),
    .X(_06812_));
 sky130_fd_sc_hd__a22o_1 _07684_ (.A1(net12),
    .A2(net35),
    .B1(net34),
    .B2(net149),
    .X(_06813_));
 sky130_fd_sc_hd__and2b_1 _07685_ (.A_N(_06812_),
    .B(_06813_),
    .X(_06814_));
 sky130_fd_sc_hd__nand2_1 _07686_ (.A(net26),
    .B(net64),
    .Y(_06815_));
 sky130_fd_sc_hd__xnor2_1 _07687_ (.A(_06814_),
    .B(_06815_),
    .Y(_06816_));
 sky130_fd_sc_hd__a31o_1 _07688_ (.A1(_01120_),
    .A2(_03499_),
    .A3(_06813_),
    .B1(_06812_),
    .X(_06817_));
 sky130_fd_sc_hd__clkbuf_4 _07689_ (.A(net35),
    .X(_06818_));
 sky130_fd_sc_hd__clkbuf_4 _07690_ (.A(_06818_),
    .X(_06819_));
 sky130_fd_sc_hd__clkbuf_4 _07691_ (.A(net34),
    .X(_06820_));
 sky130_fd_sc_hd__clkbuf_4 _07692_ (.A(_06820_),
    .X(_06821_));
 sky130_fd_sc_hd__nand4_1 _07693_ (.A(_00891_),
    .B(_01120_),
    .C(_06819_),
    .D(_06821_),
    .Y(_06822_));
 sky130_fd_sc_hd__a22o_1 _07694_ (.A1(_01076_),
    .A2(_06818_),
    .B1(_06820_),
    .B2(_01120_),
    .X(_06823_));
 sky130_fd_sc_hd__and3_2 _07695_ (.A(_06817_),
    .B(_06822_),
    .C(_06823_),
    .X(_06824_));
 sky130_fd_sc_hd__a21oi_1 _07696_ (.A1(_06822_),
    .A2(_06823_),
    .B1(_06817_),
    .Y(_06825_));
 sky130_fd_sc_hd__nor2_1 _07697_ (.A(_06824_),
    .B(_06825_),
    .Y(_06826_));
 sky130_fd_sc_hd__and3_1 _07698_ (.A(_06809_),
    .B(_06816_),
    .C(_06826_),
    .X(_06827_));
 sky130_fd_sc_hd__a21oi_1 _07699_ (.A1(_06809_),
    .A2(_06816_),
    .B1(_06826_),
    .Y(_06828_));
 sky130_fd_sc_hd__nor2_1 _07700_ (.A(_06827_),
    .B(_06828_),
    .Y(_06829_));
 sky130_fd_sc_hd__a22o_1 _07701_ (.A1(net12),
    .A2(net64),
    .B1(net34),
    .B2(net1),
    .X(_06830_));
 sky130_fd_sc_hd__and4_1 _07702_ (.A(net1),
    .B(net12),
    .C(net64),
    .D(net34),
    .X(_06831_));
 sky130_fd_sc_hd__a31o_1 _07703_ (.A1(net149),
    .A2(net63),
    .A3(_06830_),
    .B1(_06831_),
    .X(_06832_));
 sky130_fd_sc_hd__and3_1 _07704_ (.A(_01230_),
    .B(_00475_),
    .C(_06832_),
    .X(_06833_));
 sky130_fd_sc_hd__or2b_1 _07705_ (.A(_06802_),
    .B_N(_06797_),
    .X(_06834_));
 sky130_fd_sc_hd__nand2_1 _07706_ (.A(_00880_),
    .B(net64),
    .Y(_06835_));
 sky130_fd_sc_hd__xnor2_1 _07707_ (.A(_06834_),
    .B(_06835_),
    .Y(_06836_));
 sky130_fd_sc_hd__nand2_1 _07708_ (.A(net26),
    .B(net63),
    .Y(_06837_));
 sky130_fd_sc_hd__xnor2_1 _07709_ (.A(_06832_),
    .B(_06837_),
    .Y(_06838_));
 sky130_fd_sc_hd__and2b_1 _07710_ (.A_N(_06836_),
    .B(_06838_),
    .X(_06839_));
 sky130_fd_sc_hd__xor2_1 _07711_ (.A(_06809_),
    .B(_06816_),
    .X(_06840_));
 sky130_fd_sc_hd__or3_1 _07712_ (.A(_06833_),
    .B(_06839_),
    .C(_06840_),
    .X(_06841_));
 sky130_fd_sc_hd__nand2_1 _07713_ (.A(_00880_),
    .B(net63),
    .Y(_06842_));
 sky130_fd_sc_hd__and2b_1 _07714_ (.A_N(_06831_),
    .B(_06830_),
    .X(_06843_));
 sky130_fd_sc_hd__xnor2_1 _07715_ (.A(_06842_),
    .B(_06843_),
    .Y(_06844_));
 sky130_fd_sc_hd__and2_1 _07716_ (.A(_03598_),
    .B(_06844_),
    .X(_06845_));
 sky130_fd_sc_hd__xnor2_1 _07717_ (.A(_06836_),
    .B(_06838_),
    .Y(_06846_));
 sky130_fd_sc_hd__and2_1 _07718_ (.A(_06845_),
    .B(_06846_),
    .X(_06847_));
 sky130_fd_sc_hd__o21a_1 _07719_ (.A1(_06833_),
    .A2(_06839_),
    .B1(_06840_),
    .X(_06848_));
 sky130_fd_sc_hd__a21o_1 _07720_ (.A1(_06841_),
    .A2(_06847_),
    .B1(_06848_),
    .X(_06849_));
 sky130_fd_sc_hd__xor2_2 _07721_ (.A(_06829_),
    .B(_06849_),
    .X(_06850_));
 sky130_fd_sc_hd__nor2_1 _07722_ (.A(_06790_),
    .B(_06850_),
    .Y(_06851_));
 sky130_fd_sc_hd__and4_1 _07723_ (.A(_02105_),
    .B(_00650_),
    .C(_03510_),
    .D(_00475_),
    .X(_06852_));
 sky130_fd_sc_hd__a22oi_1 _07724_ (.A1(_02259_),
    .A2(_03543_),
    .B1(_00508_),
    .B2(_02171_),
    .Y(_06853_));
 sky130_fd_sc_hd__or2_1 _07725_ (.A(_06852_),
    .B(_06853_),
    .X(_06854_));
 sky130_fd_sc_hd__nand2_1 _07726_ (.A(_06790_),
    .B(_06850_),
    .Y(_06855_));
 sky130_fd_sc_hd__o21ai_1 _07727_ (.A1(_06851_),
    .A2(_06854_),
    .B1(_06855_),
    .Y(_06856_));
 sky130_fd_sc_hd__and4_1 _07728_ (.A(_00563_),
    .B(net28),
    .C(net64),
    .D(net34),
    .X(_06857_));
 sky130_fd_sc_hd__a22o_1 _07729_ (.A1(net28),
    .A2(net64),
    .B1(_06820_),
    .B2(_00563_),
    .X(_06858_));
 sky130_fd_sc_hd__and2b_1 _07730_ (.A_N(_06857_),
    .B(_06858_),
    .X(_06859_));
 sky130_fd_sc_hd__nand2_1 _07731_ (.A(_02664_),
    .B(_00475_),
    .Y(_06860_));
 sky130_fd_sc_hd__xnor2_1 _07732_ (.A(_06859_),
    .B(_06860_),
    .Y(_06861_));
 sky130_fd_sc_hd__nand2_1 _07733_ (.A(_06852_),
    .B(_06861_),
    .Y(_06862_));
 sky130_fd_sc_hd__or2_1 _07734_ (.A(_06852_),
    .B(_06861_),
    .X(_06863_));
 sky130_fd_sc_hd__and2_1 _07735_ (.A(_06862_),
    .B(_06863_),
    .X(_06864_));
 sky130_fd_sc_hd__and4_1 _07736_ (.A(_00420_),
    .B(net177),
    .C(net38),
    .D(net37),
    .X(_06865_));
 sky130_fd_sc_hd__a22o_1 _07737_ (.A1(_00420_),
    .A2(net38),
    .B1(net37),
    .B2(net177),
    .X(_06866_));
 sky130_fd_sc_hd__and2b_1 _07738_ (.A_N(_06865_),
    .B(_06866_),
    .X(_06867_));
 sky130_fd_sc_hd__nand2_1 _07739_ (.A(_01284_),
    .B(_06744_),
    .Y(_06868_));
 sky130_fd_sc_hd__xnor2_1 _07740_ (.A(_06867_),
    .B(_06868_),
    .Y(_06869_));
 sky130_fd_sc_hd__nand2_1 _07741_ (.A(_06755_),
    .B(_06869_),
    .Y(_06870_));
 sky130_fd_sc_hd__or2_1 _07742_ (.A(_06755_),
    .B(_06869_),
    .X(_06871_));
 sky130_fd_sc_hd__and2_1 _07743_ (.A(_06870_),
    .B(_06871_),
    .X(_06872_));
 sky130_fd_sc_hd__clkbuf_4 _07744_ (.A(_06819_),
    .X(_06873_));
 sky130_fd_sc_hd__clkbuf_4 _07745_ (.A(_06821_),
    .X(_06874_));
 sky130_fd_sc_hd__clkbuf_4 _07746_ (.A(_06874_),
    .X(_06875_));
 sky130_fd_sc_hd__nand2_1 _07747_ (.A(_01383_),
    .B(_06875_),
    .Y(_06876_));
 sky130_fd_sc_hd__and3_1 _07748_ (.A(_01350_),
    .B(_06873_),
    .C(_06876_),
    .X(_06877_));
 sky130_fd_sc_hd__xor2_2 _07749_ (.A(_06824_),
    .B(_06877_),
    .X(_06878_));
 sky130_fd_sc_hd__a21oi_2 _07750_ (.A1(_06829_),
    .A2(_06849_),
    .B1(_06827_),
    .Y(_06879_));
 sky130_fd_sc_hd__xnor2_2 _07751_ (.A(_06878_),
    .B(_06879_),
    .Y(_06880_));
 sky130_fd_sc_hd__xnor2_1 _07752_ (.A(_06872_),
    .B(_06880_),
    .Y(_06881_));
 sky130_fd_sc_hd__xnor2_1 _07753_ (.A(_06864_),
    .B(_06881_),
    .Y(_06882_));
 sky130_fd_sc_hd__xnor2_1 _07754_ (.A(_06856_),
    .B(_06882_),
    .Y(_06883_));
 sky130_fd_sc_hd__nand2_2 _07755_ (.A(_02259_),
    .B(_00508_),
    .Y(_06884_));
 sky130_fd_sc_hd__buf_4 _07756_ (.A(_06775_),
    .X(_06885_));
 sky130_fd_sc_hd__or2b_1 _07757_ (.A(_06848_),
    .B_N(_06841_),
    .X(_06886_));
 sky130_fd_sc_hd__xnor2_1 _07758_ (.A(_06886_),
    .B(_06847_),
    .Y(_06887_));
 sky130_fd_sc_hd__nand3_1 _07759_ (.A(_00453_),
    .B(_06885_),
    .C(_06887_),
    .Y(_06888_));
 sky130_fd_sc_hd__a21o_1 _07760_ (.A1(_00442_),
    .A2(_06775_),
    .B1(_06887_),
    .X(_06889_));
 sky130_fd_sc_hd__a21bo_1 _07761_ (.A1(_06884_),
    .A2(_06888_),
    .B1_N(_06889_),
    .X(_06890_));
 sky130_fd_sc_hd__xnor2_1 _07762_ (.A(_06790_),
    .B(_06850_),
    .Y(_06891_));
 sky130_fd_sc_hd__xnor2_1 _07763_ (.A(_06854_),
    .B(_06891_),
    .Y(_06892_));
 sky130_fd_sc_hd__nor2_1 _07764_ (.A(_06890_),
    .B(_06892_),
    .Y(_06893_));
 sky130_fd_sc_hd__xnor2_1 _07765_ (.A(_06883_),
    .B(_06893_),
    .Y(_06894_));
 sky130_fd_sc_hd__a211o_1 _07766_ (.A1(net150),
    .A2(_06175_),
    .B1(_06406_),
    .C1(_06615_),
    .X(_06895_));
 sky130_fd_sc_hd__nand3_1 _07767_ (.A(_06680_),
    .B(_06701_),
    .C(_06895_),
    .Y(_06896_));
 sky130_fd_sc_hd__and3_1 _07768_ (.A(_06723_),
    .B(_06894_),
    .C(_06896_),
    .X(_06897_));
 sky130_fd_sc_hd__a21oi_1 _07769_ (.A1(_06723_),
    .A2(_06896_),
    .B1(_06894_),
    .Y(_06898_));
 sky130_fd_sc_hd__o21bai_2 _07770_ (.A1(_05412_),
    .A2(_06897_),
    .B1_N(_06898_),
    .Y(_06899_));
 sky130_fd_sc_hd__and4_1 _07771_ (.A(_00705_),
    .B(_00573_),
    .C(_04851_),
    .D(net4),
    .X(_06900_));
 sky130_fd_sc_hd__a22o_1 _07772_ (.A1(_01208_),
    .A2(_04851_),
    .B1(net4),
    .B2(_00705_),
    .X(_06901_));
 sky130_fd_sc_hd__and2b_1 _07773_ (.A_N(_06900_),
    .B(_06901_),
    .X(_06902_));
 sky130_fd_sc_hd__nand2_1 _07774_ (.A(_01470_),
    .B(net6),
    .Y(_06903_));
 sky130_fd_sc_hd__xnor2_1 _07775_ (.A(_06902_),
    .B(_06903_),
    .Y(_06904_));
 sky130_fd_sc_hd__a31o_1 _07776_ (.A1(net33),
    .A2(net6),
    .A3(_05005_),
    .B1(_04994_),
    .X(_06905_));
 sky130_fd_sc_hd__and2_1 _07777_ (.A(net33),
    .B(net7),
    .X(_06906_));
 sky130_fd_sc_hd__xor2_1 _07778_ (.A(_06905_),
    .B(_06906_),
    .X(_06907_));
 sky130_fd_sc_hd__xnor2_1 _07779_ (.A(_06904_),
    .B(_06907_),
    .Y(_06908_));
 sky130_fd_sc_hd__nor2_1 _07780_ (.A(_05060_),
    .B(_06908_),
    .Y(_06909_));
 sky130_fd_sc_hd__and2_1 _07781_ (.A(_05060_),
    .B(_06908_),
    .X(_06910_));
 sky130_fd_sc_hd__or2_1 _07782_ (.A(_06909_),
    .B(_06910_),
    .X(_06911_));
 sky130_fd_sc_hd__and4_1 _07783_ (.A(_01044_),
    .B(_03147_),
    .C(_00355_),
    .D(_02960_),
    .X(_06912_));
 sky130_fd_sc_hd__a22o_1 _07784_ (.A1(_01044_),
    .A2(_00355_),
    .B1(_02960_),
    .B2(_03147_),
    .X(_06913_));
 sky130_fd_sc_hd__and2b_1 _07785_ (.A_N(_06912_),
    .B(_06913_),
    .X(_06914_));
 sky130_fd_sc_hd__nand2_1 _07786_ (.A(_01000_),
    .B(_04378_),
    .Y(_06915_));
 sky130_fd_sc_hd__xnor2_1 _07787_ (.A(_06914_),
    .B(_06915_),
    .Y(_06916_));
 sky130_fd_sc_hd__a31o_1 _07788_ (.A1(net59),
    .A2(_04367_),
    .A3(_05104_),
    .B1(_05093_),
    .X(_06917_));
 sky130_fd_sc_hd__nand2_1 _07789_ (.A(net59),
    .B(_04455_),
    .Y(_06918_));
 sky130_fd_sc_hd__xnor2_1 _07790_ (.A(_06917_),
    .B(_06918_),
    .Y(_06919_));
 sky130_fd_sc_hd__xnor2_1 _07791_ (.A(_06916_),
    .B(_06919_),
    .Y(_06920_));
 sky130_fd_sc_hd__nor2_2 _07792_ (.A(_05148_),
    .B(_06920_),
    .Y(_06921_));
 sky130_fd_sc_hd__and2_1 _07793_ (.A(_05148_),
    .B(_06920_),
    .X(_06922_));
 sky130_fd_sc_hd__nor2_1 _07794_ (.A(_06921_),
    .B(_06922_),
    .Y(_06923_));
 sky130_fd_sc_hd__and2b_1 _07795_ (.A_N(_05236_),
    .B(_05258_),
    .X(_06924_));
 sky130_fd_sc_hd__a21bo_1 _07796_ (.A1(_04532_),
    .A2(_05225_),
    .B1_N(_04499_),
    .X(_06925_));
 sky130_fd_sc_hd__or3_4 _07797_ (.A(_06923_),
    .B(_06924_),
    .C(_06925_),
    .X(_06926_));
 sky130_fd_sc_hd__o21ai_1 _07798_ (.A1(_06924_),
    .A2(_06925_),
    .B1(_06923_),
    .Y(_06927_));
 sky130_fd_sc_hd__nand2_2 _07799_ (.A(_06926_),
    .B(_06927_),
    .Y(_06928_));
 sky130_fd_sc_hd__xor2_2 _07800_ (.A(_06911_),
    .B(_06928_),
    .X(_06929_));
 sky130_fd_sc_hd__o21ba_1 _07801_ (.A1(_05170_),
    .A2(_05269_),
    .B1_N(_05082_),
    .X(_06930_));
 sky130_fd_sc_hd__a21o_1 _07802_ (.A1(_05170_),
    .A2(_05269_),
    .B1(_06930_),
    .X(_06931_));
 sky130_fd_sc_hd__xnor2_1 _07803_ (.A(_06929_),
    .B(_06931_),
    .Y(_06932_));
 sky130_fd_sc_hd__nand2_1 _07804_ (.A(_04983_),
    .B(_05291_),
    .Y(_06933_));
 sky130_fd_sc_hd__o31ai_2 _07805_ (.A1(_05302_),
    .A2(_05368_),
    .A3(_05390_),
    .B1(_06933_),
    .Y(_06934_));
 sky130_fd_sc_hd__xnor2_2 _07806_ (.A(net148),
    .B(net166),
    .Y(_06935_));
 sky130_fd_sc_hd__and2_1 _07807_ (.A(_06658_),
    .B(_06669_),
    .X(_06936_));
 sky130_fd_sc_hd__buf_4 _07808_ (.A(_06472_),
    .X(_06937_));
 sky130_fd_sc_hd__and4_1 _07809_ (.A(_06626_),
    .B(_06450_),
    .C(_06937_),
    .D(_06637_),
    .X(_06938_));
 sky130_fd_sc_hd__a211o_1 _07810_ (.A1(_06527_),
    .A2(_06648_),
    .B1(_06936_),
    .C1(_06938_),
    .X(_06939_));
 sky130_fd_sc_hd__and4_1 _07811_ (.A(net27),
    .B(net28),
    .C(_06818_),
    .D(net34),
    .X(_06940_));
 sky130_fd_sc_hd__a22o_1 _07812_ (.A1(_00563_),
    .A2(_06818_),
    .B1(_06820_),
    .B2(_00639_),
    .X(_06941_));
 sky130_fd_sc_hd__and2b_1 _07813_ (.A_N(_06940_),
    .B(_06941_),
    .X(_06942_));
 sky130_fd_sc_hd__nand2_1 _07814_ (.A(_00541_),
    .B(_03499_),
    .Y(_06943_));
 sky130_fd_sc_hd__xnor2_1 _07815_ (.A(_06942_),
    .B(_06943_),
    .Y(_06944_));
 sky130_fd_sc_hd__a31o_1 _07816_ (.A1(net29),
    .A2(net63),
    .A3(_06858_),
    .B1(_06857_),
    .X(_06945_));
 sky130_fd_sc_hd__nand2_1 _07817_ (.A(_02719_),
    .B(net63),
    .Y(_06946_));
 sky130_fd_sc_hd__xnor2_1 _07818_ (.A(_06945_),
    .B(_06946_),
    .Y(_06947_));
 sky130_fd_sc_hd__xnor2_1 _07819_ (.A(_06944_),
    .B(_06947_),
    .Y(_06948_));
 sky130_fd_sc_hd__nor2_1 _07820_ (.A(_06862_),
    .B(_06948_),
    .Y(_06949_));
 sky130_fd_sc_hd__and2_1 _07821_ (.A(_06862_),
    .B(_06948_),
    .X(_06950_));
 sky130_fd_sc_hd__or2_1 _07822_ (.A(_06949_),
    .B(_06950_),
    .X(_06951_));
 sky130_fd_sc_hd__and4_1 _07823_ (.A(_00420_),
    .B(net177),
    .C(net39),
    .D(net38),
    .X(_06952_));
 sky130_fd_sc_hd__a22o_1 _07824_ (.A1(_00420_),
    .A2(net39),
    .B1(net38),
    .B2(net177),
    .X(_06953_));
 sky130_fd_sc_hd__and2b_1 _07825_ (.A_N(_06952_),
    .B(_06953_),
    .X(_06954_));
 sky130_fd_sc_hd__nand2_1 _07826_ (.A(_01076_),
    .B(net37),
    .Y(_06955_));
 sky130_fd_sc_hd__xnor2_1 _07827_ (.A(_06954_),
    .B(_06955_),
    .Y(_06956_));
 sky130_fd_sc_hd__a31o_1 _07828_ (.A1(_00880_),
    .A2(net36),
    .A3(_06866_),
    .B1(_06865_),
    .X(_06957_));
 sky130_fd_sc_hd__nand2_1 _07829_ (.A(_01120_),
    .B(_06744_),
    .Y(_06958_));
 sky130_fd_sc_hd__xnor2_1 _07830_ (.A(_06957_),
    .B(_06958_),
    .Y(_06959_));
 sky130_fd_sc_hd__xnor2_1 _07831_ (.A(_06956_),
    .B(_06959_),
    .Y(_06960_));
 sky130_fd_sc_hd__nor2_1 _07832_ (.A(_06870_),
    .B(_06960_),
    .Y(_06961_));
 sky130_fd_sc_hd__and2_1 _07833_ (.A(_06870_),
    .B(_06960_),
    .X(_06962_));
 sky130_fd_sc_hd__nor2_1 _07834_ (.A(_06961_),
    .B(_06962_),
    .Y(_06963_));
 sky130_fd_sc_hd__clkbuf_4 _07835_ (.A(_06873_),
    .X(_06964_));
 sky130_fd_sc_hd__clkbuf_4 _07836_ (.A(_06964_),
    .X(_06965_));
 sky130_fd_sc_hd__clkbuf_4 _07837_ (.A(_06875_),
    .X(_06966_));
 sky130_fd_sc_hd__and4_1 _07838_ (.A(_01383_),
    .B(_01350_),
    .C(_06965_),
    .D(_06966_),
    .X(_06967_));
 sky130_fd_sc_hd__and2_1 _07839_ (.A(_06824_),
    .B(_06877_),
    .X(_06968_));
 sky130_fd_sc_hd__and2b_1 _07840_ (.A_N(_06878_),
    .B(_06879_),
    .X(_06969_));
 sky130_fd_sc_hd__or4_1 _07841_ (.A(_06963_),
    .B(_06967_),
    .C(_06968_),
    .D(_06969_),
    .X(_06970_));
 sky130_fd_sc_hd__o31ai_1 _07842_ (.A1(_06967_),
    .A2(_06968_),
    .A3(_06969_),
    .B1(_06963_),
    .Y(_06971_));
 sky130_fd_sc_hd__nand2_1 _07843_ (.A(_06970_),
    .B(_06971_),
    .Y(_06972_));
 sky130_fd_sc_hd__xor2_1 _07844_ (.A(_06951_),
    .B(_06972_),
    .X(_06973_));
 sky130_fd_sc_hd__a21o_1 _07845_ (.A1(_06872_),
    .A2(_06880_),
    .B1(_06864_),
    .X(_06974_));
 sky130_fd_sc_hd__o21ai_1 _07846_ (.A1(_06872_),
    .A2(_06880_),
    .B1(_06974_),
    .Y(_06975_));
 sky130_fd_sc_hd__xnor2_1 _07847_ (.A(_06973_),
    .B(_06975_),
    .Y(_06976_));
 sky130_fd_sc_hd__inv_2 _07848_ (.A(_06893_),
    .Y(_06977_));
 sky130_fd_sc_hd__nand2_1 _07849_ (.A(_06856_),
    .B(_06882_),
    .Y(_06978_));
 sky130_fd_sc_hd__o21ai_1 _07850_ (.A1(_06883_),
    .A2(_06977_),
    .B1(_06978_),
    .Y(_06979_));
 sky130_fd_sc_hd__xor2_1 _07851_ (.A(_06976_),
    .B(_06979_),
    .X(_06980_));
 sky130_fd_sc_hd__or4_4 _07852_ (.A(net139),
    .B(_06712_),
    .C(_06939_),
    .D(_06980_),
    .X(_06981_));
 sky130_fd_sc_hd__o31ai_2 _07853_ (.A1(net139),
    .A2(_06712_),
    .A3(_06939_),
    .B1(_06980_),
    .Y(_06982_));
 sky130_fd_sc_hd__nand2_2 _07854_ (.A(_06981_),
    .B(_06982_),
    .Y(_06983_));
 sky130_fd_sc_hd__xor2_2 _07855_ (.A(_06935_),
    .B(_06983_),
    .X(_06984_));
 sky130_fd_sc_hd__and2b_1 _07856_ (.A_N(_06899_),
    .B(_06984_),
    .X(_06985_));
 sky130_fd_sc_hd__or3_4 _07857_ (.A(_06898_),
    .B(_05412_),
    .C(_06897_),
    .X(_06986_));
 sky130_fd_sc_hd__o21ai_1 _07858_ (.A1(_06898_),
    .A2(_06897_),
    .B1(_05412_),
    .Y(_06987_));
 sky130_fd_sc_hd__and2_1 _07859_ (.A(_05368_),
    .B(_05390_),
    .X(_06988_));
 sky130_fd_sc_hd__nor2_1 _07860_ (.A(_05401_),
    .B(_06988_),
    .Y(_06989_));
 sky130_fd_sc_hd__a21oi_1 _07861_ (.A1(_06142_),
    .A2(_06175_),
    .B1(_06406_),
    .Y(_06990_));
 sky130_fd_sc_hd__or3_1 _07862_ (.A(_06384_),
    .B(_06615_),
    .C(_06990_),
    .X(_06991_));
 sky130_fd_sc_hd__o21ai_1 _07863_ (.A1(_06384_),
    .A2(_06990_),
    .B1(_06615_),
    .Y(_06992_));
 sky130_fd_sc_hd__nand2_1 _07864_ (.A(_06890_),
    .B(_06892_),
    .Y(_06993_));
 sky130_fd_sc_hd__nand2_1 _07865_ (.A(_06977_),
    .B(_06993_),
    .Y(_06994_));
 sky130_fd_sc_hd__a21oi_1 _07866_ (.A1(_06991_),
    .A2(_06992_),
    .B1(_06994_),
    .Y(_06995_));
 sky130_fd_sc_hd__and3_1 _07867_ (.A(_06994_),
    .B(_06991_),
    .C(_06992_),
    .X(_06996_));
 sky130_fd_sc_hd__o21bai_1 _07868_ (.A1(_06989_),
    .A2(_06995_),
    .B1_N(_06996_),
    .Y(_06997_));
 sky130_fd_sc_hd__a21o_4 _07869_ (.A1(_06986_),
    .A2(_06987_),
    .B1(_06997_),
    .X(_06998_));
 sky130_fd_sc_hd__xor2_2 _07870_ (.A(_06984_),
    .B(_06899_),
    .X(_06999_));
 sky130_fd_sc_hd__nor2_1 _07871_ (.A(_06998_),
    .B(_06999_),
    .Y(_07000_));
 sky130_fd_sc_hd__nand2_1 _07872_ (.A(_00530_),
    .B(_00410_),
    .Y(_07001_));
 sky130_fd_sc_hd__and2b_1 _07873_ (.A_N(_06975_),
    .B(_06973_),
    .X(_07002_));
 sky130_fd_sc_hd__a21o_1 _07874_ (.A1(_06976_),
    .A2(_06979_),
    .B1(_07002_),
    .X(_07003_));
 sky130_fd_sc_hd__buf_4 _07875_ (.A(_06885_),
    .X(_07004_));
 sky130_fd_sc_hd__nand2_1 _07876_ (.A(_02467_),
    .B(_07004_),
    .Y(_07005_));
 sky130_fd_sc_hd__nand2_1 _07877_ (.A(_06951_),
    .B(_06971_),
    .Y(_07006_));
 sky130_fd_sc_hd__and3_1 _07878_ (.A(_01230_),
    .B(_06744_),
    .C(_06957_),
    .X(_07007_));
 sky130_fd_sc_hd__a21o_1 _07879_ (.A1(_06956_),
    .A2(_06959_),
    .B1(_07007_),
    .X(_07008_));
 sky130_fd_sc_hd__a31o_1 _07880_ (.A1(_00891_),
    .A2(net37),
    .A3(_06953_),
    .B1(_06952_),
    .X(_07009_));
 sky130_fd_sc_hd__clkbuf_4 _07881_ (.A(net39),
    .X(_07010_));
 sky130_fd_sc_hd__a22oi_1 _07882_ (.A1(_00978_),
    .A2(_07010_),
    .B1(net38),
    .B2(net149),
    .Y(_07011_));
 sky130_fd_sc_hd__and4_1 _07883_ (.A(net177),
    .B(net149),
    .C(net39),
    .D(net38),
    .X(_07012_));
 sky130_fd_sc_hd__nor2_1 _07884_ (.A(_07011_),
    .B(_07012_),
    .Y(_07013_));
 sky130_fd_sc_hd__nand2_1 _07885_ (.A(_01120_),
    .B(net37),
    .Y(_07014_));
 sky130_fd_sc_hd__xnor2_1 _07886_ (.A(_07013_),
    .B(_07014_),
    .Y(_07015_));
 sky130_fd_sc_hd__xor2_1 _07887_ (.A(_07009_),
    .B(_07015_),
    .X(_07016_));
 sky130_fd_sc_hd__xor2_1 _07888_ (.A(_07008_),
    .B(_07016_),
    .X(_07017_));
 sky130_fd_sc_hd__xnor2_1 _07889_ (.A(_06961_),
    .B(_07017_),
    .Y(_07018_));
 sky130_fd_sc_hd__and3_1 _07890_ (.A(_02719_),
    .B(_00475_),
    .C(_06945_),
    .X(_07019_));
 sky130_fd_sc_hd__a21o_1 _07891_ (.A1(_06944_),
    .A2(_06947_),
    .B1(_07019_),
    .X(_07020_));
 sky130_fd_sc_hd__a31o_1 _07892_ (.A1(_00541_),
    .A2(_03499_),
    .A3(_06941_),
    .B1(_06940_),
    .X(_07021_));
 sky130_fd_sc_hd__a22oi_1 _07893_ (.A1(_00639_),
    .A2(_06818_),
    .B1(_06820_),
    .B2(net29),
    .Y(_07022_));
 sky130_fd_sc_hd__and4_1 _07894_ (.A(net28),
    .B(net29),
    .C(_06818_),
    .D(net34),
    .X(_07023_));
 sky130_fd_sc_hd__nor2_1 _07895_ (.A(_07022_),
    .B(_07023_),
    .Y(_07024_));
 sky130_fd_sc_hd__nand2_1 _07896_ (.A(_02719_),
    .B(_03499_),
    .Y(_07025_));
 sky130_fd_sc_hd__xnor2_1 _07897_ (.A(_07024_),
    .B(_07025_),
    .Y(_07026_));
 sky130_fd_sc_hd__xor2_1 _07898_ (.A(_07021_),
    .B(_07026_),
    .X(_07027_));
 sky130_fd_sc_hd__xor2_1 _07899_ (.A(_07020_),
    .B(_07027_),
    .X(_07028_));
 sky130_fd_sc_hd__xnor2_1 _07900_ (.A(_06949_),
    .B(_07028_),
    .Y(_07029_));
 sky130_fd_sc_hd__nor2_1 _07901_ (.A(_07018_),
    .B(_07029_),
    .Y(_07030_));
 sky130_fd_sc_hd__and2_1 _07902_ (.A(_07018_),
    .B(_07029_),
    .X(_07031_));
 sky130_fd_sc_hd__nor2_1 _07903_ (.A(_07030_),
    .B(_07031_),
    .Y(_07032_));
 sky130_fd_sc_hd__a21oi_1 _07904_ (.A1(_06970_),
    .A2(_07006_),
    .B1(_07032_),
    .Y(_07033_));
 sky130_fd_sc_hd__nand3_1 _07905_ (.A(_06970_),
    .B(_07032_),
    .C(_07006_),
    .Y(_07034_));
 sky130_fd_sc_hd__or2b_1 _07906_ (.A(_07033_),
    .B_N(_07034_),
    .X(_07035_));
 sky130_fd_sc_hd__xor2_2 _07907_ (.A(_07005_),
    .B(_07035_),
    .X(_07036_));
 sky130_fd_sc_hd__xor2_1 _07908_ (.A(_07003_),
    .B(_07036_),
    .X(_07037_));
 sky130_fd_sc_hd__and2b_1 _07909_ (.A_N(_06931_),
    .B(_06929_),
    .X(_07038_));
 sky130_fd_sc_hd__a21o_1 _07910_ (.A1(_06932_),
    .A2(_06934_),
    .B1(_07038_),
    .X(_07039_));
 sky130_fd_sc_hd__buf_4 _07911_ (.A(_04939_),
    .X(_07040_));
 sky130_fd_sc_hd__nand2_2 _07912_ (.A(_02456_),
    .B(_07040_),
    .Y(_07041_));
 sky130_fd_sc_hd__nand2_1 _07913_ (.A(_06911_),
    .B(_06927_),
    .Y(_07042_));
 sky130_fd_sc_hd__and3_1 _07914_ (.A(_00901_),
    .B(_04455_),
    .C(_06917_),
    .X(_07043_));
 sky130_fd_sc_hd__a21o_1 _07915_ (.A1(_06916_),
    .A2(_06919_),
    .B1(_07043_),
    .X(_07044_));
 sky130_fd_sc_hd__a31o_1 _07916_ (.A1(_01996_),
    .A2(_04378_),
    .A3(_06913_),
    .B1(_06912_),
    .X(_07045_));
 sky130_fd_sc_hd__a22oi_1 _07917_ (.A1(net62),
    .A2(net32),
    .B1(_04367_),
    .B2(net61),
    .Y(_07046_));
 sky130_fd_sc_hd__and4_1 _07918_ (.A(net62),
    .B(net61),
    .C(net32),
    .D(net2),
    .X(_07047_));
 sky130_fd_sc_hd__and4bb_1 _07919_ (.A_N(_07046_),
    .B_N(_07047_),
    .C(net60),
    .D(net3),
    .X(_07048_));
 sky130_fd_sc_hd__o2bb2a_1 _07920_ (.A1_N(_01000_),
    .A2_N(_04455_),
    .B1(_07046_),
    .B2(net173),
    .X(_07049_));
 sky130_fd_sc_hd__nor2_1 _07921_ (.A(_07048_),
    .B(_07049_),
    .Y(_07050_));
 sky130_fd_sc_hd__xor2_1 _07922_ (.A(_07045_),
    .B(_07050_),
    .X(_07051_));
 sky130_fd_sc_hd__and2_1 _07923_ (.A(_07044_),
    .B(_07051_),
    .X(_07052_));
 sky130_fd_sc_hd__or2_1 _07924_ (.A(_07044_),
    .B(_07051_),
    .X(_07053_));
 sky130_fd_sc_hd__and2b_1 _07925_ (.A_N(_07052_),
    .B(_07053_),
    .X(_07054_));
 sky130_fd_sc_hd__xnor2_1 _07926_ (.A(_06921_),
    .B(_07054_),
    .Y(_07055_));
 sky130_fd_sc_hd__nand2_1 _07927_ (.A(_06905_),
    .B(_06906_),
    .Y(_07056_));
 sky130_fd_sc_hd__a21bo_1 _07928_ (.A1(_06904_),
    .A2(_06907_),
    .B1_N(_07056_),
    .X(_07057_));
 sky130_fd_sc_hd__a31o_1 _07929_ (.A1(_00672_),
    .A2(_05027_),
    .A3(_06901_),
    .B1(_06900_),
    .X(_07058_));
 sky130_fd_sc_hd__a22oi_1 _07930_ (.A1(net163),
    .A2(net6),
    .B1(net5),
    .B2(_00705_),
    .Y(_07059_));
 sky130_fd_sc_hd__and4_1 _07931_ (.A(net58),
    .B(_00716_),
    .C(net6),
    .D(net5),
    .X(_07060_));
 sky130_fd_sc_hd__and4bb_1 _07932_ (.A_N(_07059_),
    .B_N(_07060_),
    .C(net44),
    .D(net7),
    .X(_07061_));
 sky130_fd_sc_hd__o2bb2a_1 _07933_ (.A1_N(_01470_),
    .A2_N(net7),
    .B1(_07059_),
    .B2(_07060_),
    .X(_07062_));
 sky130_fd_sc_hd__nor2_1 _07934_ (.A(net172),
    .B(_07062_),
    .Y(_07063_));
 sky130_fd_sc_hd__xor2_1 _07935_ (.A(_07058_),
    .B(_07063_),
    .X(_07064_));
 sky130_fd_sc_hd__and2_1 _07936_ (.A(_07057_),
    .B(_07064_),
    .X(_07065_));
 sky130_fd_sc_hd__or2_1 _07937_ (.A(_07057_),
    .B(_07064_),
    .X(_07066_));
 sky130_fd_sc_hd__and2b_1 _07938_ (.A_N(_07065_),
    .B(_07066_),
    .X(_07067_));
 sky130_fd_sc_hd__xnor2_1 _07939_ (.A(_06909_),
    .B(_07067_),
    .Y(_07068_));
 sky130_fd_sc_hd__nor2_1 _07940_ (.A(_07055_),
    .B(_07068_),
    .Y(_07069_));
 sky130_fd_sc_hd__and2_1 _07941_ (.A(_07055_),
    .B(_07068_),
    .X(_07070_));
 sky130_fd_sc_hd__nor2_1 _07942_ (.A(_07069_),
    .B(_07070_),
    .Y(_07071_));
 sky130_fd_sc_hd__a21oi_1 _07943_ (.A1(_06926_),
    .A2(_07042_),
    .B1(_07071_),
    .Y(_07072_));
 sky130_fd_sc_hd__nand3_1 _07944_ (.A(_06926_),
    .B(_07071_),
    .C(_07042_),
    .Y(_07073_));
 sky130_fd_sc_hd__and2b_1 _07945_ (.A_N(_07073_),
    .B(_07072_),
    .X(_07074_));
 sky130_fd_sc_hd__xnor2_4 _07946_ (.A(_07041_),
    .B(_07074_),
    .Y(_07075_));
 sky130_fd_sc_hd__xor2_1 _07947_ (.A(net165),
    .B(_07075_),
    .X(_07076_));
 sky130_fd_sc_hd__and2_1 _07948_ (.A(_07037_),
    .B(_07076_),
    .X(_07077_));
 sky130_fd_sc_hd__nor2_1 _07949_ (.A(_07037_),
    .B(_07076_),
    .Y(_07078_));
 sky130_fd_sc_hd__nor2_1 _07950_ (.A(_07077_),
    .B(_07078_),
    .Y(_07079_));
 sky130_fd_sc_hd__a21boi_4 _07951_ (.A1(_06935_),
    .A2(_06982_),
    .B1_N(_06981_),
    .Y(_07080_));
 sky130_fd_sc_hd__xor2_2 _07952_ (.A(_07079_),
    .B(_07080_),
    .X(_07081_));
 sky130_fd_sc_hd__xnor2_2 _07953_ (.A(_07001_),
    .B(_07081_),
    .Y(_07082_));
 sky130_fd_sc_hd__o21a_1 _07954_ (.A1(_06985_),
    .A2(_07000_),
    .B1(_07082_),
    .X(_07083_));
 sky130_fd_sc_hd__and4_1 _07955_ (.A(_03532_),
    .B(_00497_),
    .C(_00388_),
    .D(_03004_),
    .X(_07084_));
 sky130_fd_sc_hd__inv_2 _07956_ (.A(_07084_),
    .Y(_00000_));
 sky130_fd_sc_hd__a22o_1 _07957_ (.A1(_03554_),
    .A2(_00410_),
    .B1(_03015_),
    .B2(_00519_),
    .X(_00001_));
 sky130_fd_sc_hd__and2_1 _07958_ (.A(_00000_),
    .B(_00001_),
    .X(_00002_));
 sky130_fd_sc_hd__clkbuf_4 _07959_ (.A(_06765_),
    .X(_00003_));
 sky130_fd_sc_hd__clkbuf_4 _07960_ (.A(_00003_),
    .X(_00004_));
 sky130_fd_sc_hd__a22oi_1 _07961_ (.A1(_02259_),
    .A2(_00004_),
    .B1(_07004_),
    .B2(_02171_),
    .Y(_00005_));
 sky130_fd_sc_hd__and4_1 _07962_ (.A(_02259_),
    .B(_02171_),
    .C(_00004_),
    .D(_06885_),
    .X(_00006_));
 sky130_fd_sc_hd__nor2_1 _07963_ (.A(_00005_),
    .B(_00006_),
    .Y(_00007_));
 sky130_fd_sc_hd__nand2_1 _07964_ (.A(_07009_),
    .B(_07015_),
    .Y(_00008_));
 sky130_fd_sc_hd__a31o_1 _07965_ (.A1(_01120_),
    .A2(net37),
    .A3(_07013_),
    .B1(_07012_),
    .X(_00009_));
 sky130_fd_sc_hd__a22o_1 _07966_ (.A1(_01076_),
    .A2(_07010_),
    .B1(net38),
    .B2(_01120_),
    .X(_00010_));
 sky130_fd_sc_hd__nand4_1 _07967_ (.A(_00891_),
    .B(_01120_),
    .C(_07010_),
    .D(net38),
    .Y(_00011_));
 sky130_fd_sc_hd__nand2_1 _07968_ (.A(_00010_),
    .B(_00011_),
    .Y(_00012_));
 sky130_fd_sc_hd__xor2_1 _07969_ (.A(_00009_),
    .B(_00012_),
    .X(_00013_));
 sky130_fd_sc_hd__nor2_1 _07970_ (.A(_00008_),
    .B(_00013_),
    .Y(_00014_));
 sky130_fd_sc_hd__and2_1 _07971_ (.A(_00008_),
    .B(_00013_),
    .X(_00015_));
 sky130_fd_sc_hd__or2_1 _07972_ (.A(_00014_),
    .B(_00015_),
    .X(_00016_));
 sky130_fd_sc_hd__and2_1 _07973_ (.A(_07008_),
    .B(_07016_),
    .X(_00017_));
 sky130_fd_sc_hd__a21oi_1 _07974_ (.A1(_06961_),
    .A2(_07017_),
    .B1(_00017_),
    .Y(_00018_));
 sky130_fd_sc_hd__xor2_1 _07975_ (.A(_00016_),
    .B(_00018_),
    .X(_00019_));
 sky130_fd_sc_hd__nand2_1 _07976_ (.A(_07021_),
    .B(_07026_),
    .Y(_00020_));
 sky130_fd_sc_hd__a31o_1 _07977_ (.A1(_02719_),
    .A2(_03499_),
    .A3(_07024_),
    .B1(_07023_),
    .X(_00021_));
 sky130_fd_sc_hd__a22o_1 _07978_ (.A1(_00541_),
    .A2(_06818_),
    .B1(_06821_),
    .B2(net30),
    .X(_00022_));
 sky130_fd_sc_hd__nand4_1 _07979_ (.A(_00541_),
    .B(_02719_),
    .C(_06819_),
    .D(_06821_),
    .Y(_00023_));
 sky130_fd_sc_hd__nand2_1 _07980_ (.A(_00022_),
    .B(_00023_),
    .Y(_00024_));
 sky130_fd_sc_hd__xor2_1 _07981_ (.A(_00021_),
    .B(_00024_),
    .X(_00025_));
 sky130_fd_sc_hd__nor2_1 _07982_ (.A(_00020_),
    .B(_00025_),
    .Y(_00026_));
 sky130_fd_sc_hd__and2_1 _07983_ (.A(_00020_),
    .B(_00025_),
    .X(_00027_));
 sky130_fd_sc_hd__or2_1 _07984_ (.A(_00026_),
    .B(_00027_),
    .X(_00028_));
 sky130_fd_sc_hd__and2_1 _07985_ (.A(_07020_),
    .B(_07027_),
    .X(_00029_));
 sky130_fd_sc_hd__a21oi_1 _07986_ (.A1(_06949_),
    .A2(_07028_),
    .B1(_00029_),
    .Y(_00030_));
 sky130_fd_sc_hd__xor2_1 _07987_ (.A(_00028_),
    .B(_00030_),
    .X(_00031_));
 sky130_fd_sc_hd__nand2_1 _07988_ (.A(_00019_),
    .B(_00031_),
    .Y(_00032_));
 sky130_fd_sc_hd__or2_1 _07989_ (.A(_00019_),
    .B(_00031_),
    .X(_00033_));
 sky130_fd_sc_hd__and2_1 _07990_ (.A(_00032_),
    .B(_00033_),
    .X(_00034_));
 sky130_fd_sc_hd__nand2_1 _07991_ (.A(_07030_),
    .B(_00034_),
    .Y(_00035_));
 sky130_fd_sc_hd__or2_1 _07992_ (.A(_07030_),
    .B(_00034_),
    .X(_00036_));
 sky130_fd_sc_hd__nand2_1 _07993_ (.A(_00035_),
    .B(_00036_),
    .Y(_00037_));
 sky130_fd_sc_hd__xor2_1 _07994_ (.A(_00007_),
    .B(_00037_),
    .X(_00038_));
 sky130_fd_sc_hd__a21o_1 _07995_ (.A1(_07005_),
    .A2(_07034_),
    .B1(_07033_),
    .X(_00039_));
 sky130_fd_sc_hd__xor2_1 _07996_ (.A(_00038_),
    .B(_00039_),
    .X(_00040_));
 sky130_fd_sc_hd__and3_1 _07997_ (.A(_07003_),
    .B(_07036_),
    .C(_00040_),
    .X(_00041_));
 sky130_fd_sc_hd__a21oi_1 _07998_ (.A1(_07003_),
    .A2(_07036_),
    .B1(_00040_),
    .Y(_00042_));
 sky130_fd_sc_hd__a22o_1 _07999_ (.A1(_02335_),
    .A2(_04917_),
    .B1(_04939_),
    .B2(_03070_),
    .X(_00043_));
 sky130_fd_sc_hd__and4_1 _08000_ (.A(_03059_),
    .B(_02040_),
    .C(_04917_),
    .D(_04939_),
    .X(_00044_));
 sky130_fd_sc_hd__inv_2 _08001_ (.A(_00044_),
    .Y(_00045_));
 sky130_fd_sc_hd__and2_1 _08002_ (.A(_00043_),
    .B(_00045_),
    .X(_00046_));
 sky130_fd_sc_hd__nand2_1 _08003_ (.A(_07045_),
    .B(_07050_),
    .Y(_00047_));
 sky130_fd_sc_hd__a22o_1 _08004_ (.A1(_01044_),
    .A2(_04367_),
    .B1(net3),
    .B2(_03147_),
    .X(_00048_));
 sky130_fd_sc_hd__nand4_1 _08005_ (.A(_01044_),
    .B(_03147_),
    .C(_04367_),
    .D(_04455_),
    .Y(_00049_));
 sky130_fd_sc_hd__o211a_1 _08006_ (.A1(_07047_),
    .A2(_07048_),
    .B1(_00048_),
    .C1(_00049_),
    .X(_00050_));
 sky130_fd_sc_hd__a211oi_1 _08007_ (.A1(_00048_),
    .A2(_00049_),
    .B1(net174),
    .C1(_07048_),
    .Y(_00051_));
 sky130_fd_sc_hd__or2_1 _08008_ (.A(_00050_),
    .B(_00051_),
    .X(_00052_));
 sky130_fd_sc_hd__nor2_1 _08009_ (.A(_00047_),
    .B(_00052_),
    .Y(_00053_));
 sky130_fd_sc_hd__and2_1 _08010_ (.A(_00047_),
    .B(_00052_),
    .X(_00054_));
 sky130_fd_sc_hd__or2_1 _08011_ (.A(_00053_),
    .B(_00054_),
    .X(_00055_));
 sky130_fd_sc_hd__a21oi_1 _08012_ (.A1(_06921_),
    .A2(_07053_),
    .B1(_07052_),
    .Y(_00056_));
 sky130_fd_sc_hd__xor2_1 _08013_ (.A(_00055_),
    .B(_00056_),
    .X(_00057_));
 sky130_fd_sc_hd__nand2_1 _08014_ (.A(_07058_),
    .B(_07063_),
    .Y(_00058_));
 sky130_fd_sc_hd__a22o_1 _08015_ (.A1(_01197_),
    .A2(net6),
    .B1(net7),
    .B2(_01208_),
    .X(_00059_));
 sky130_fd_sc_hd__nand4_1 _08016_ (.A(_01197_),
    .B(_04510_),
    .C(net6),
    .D(net7),
    .Y(_00060_));
 sky130_fd_sc_hd__o211a_1 _08017_ (.A1(net159),
    .A2(_07061_),
    .B1(_00059_),
    .C1(_00060_),
    .X(_00061_));
 sky130_fd_sc_hd__a211oi_1 _08018_ (.A1(_00059_),
    .A2(_00060_),
    .B1(net158),
    .C1(net171),
    .Y(_00062_));
 sky130_fd_sc_hd__or2_1 _08019_ (.A(_00061_),
    .B(_00062_),
    .X(_00063_));
 sky130_fd_sc_hd__nor2_1 _08020_ (.A(_00058_),
    .B(_00063_),
    .Y(_00064_));
 sky130_fd_sc_hd__and2_1 _08021_ (.A(_00058_),
    .B(_00063_),
    .X(_00065_));
 sky130_fd_sc_hd__or2_1 _08022_ (.A(_00064_),
    .B(_00065_),
    .X(_00066_));
 sky130_fd_sc_hd__a21oi_1 _08023_ (.A1(_06909_),
    .A2(_07066_),
    .B1(_07065_),
    .Y(_00067_));
 sky130_fd_sc_hd__xor2_1 _08024_ (.A(_00066_),
    .B(_00067_),
    .X(_00068_));
 sky130_fd_sc_hd__nand2_1 _08025_ (.A(_00057_),
    .B(_00068_),
    .Y(_00069_));
 sky130_fd_sc_hd__or2_1 _08026_ (.A(_00057_),
    .B(_00068_),
    .X(_00070_));
 sky130_fd_sc_hd__and2_1 _08027_ (.A(_00069_),
    .B(_00070_),
    .X(_00071_));
 sky130_fd_sc_hd__nand2_1 _08028_ (.A(_07069_),
    .B(_00071_),
    .Y(_00072_));
 sky130_fd_sc_hd__or2_1 _08029_ (.A(_07069_),
    .B(_00071_),
    .X(_00073_));
 sky130_fd_sc_hd__nand2_1 _08030_ (.A(_00072_),
    .B(_00073_),
    .Y(_00074_));
 sky130_fd_sc_hd__xor2_2 _08031_ (.A(_00046_),
    .B(_00074_),
    .X(_00075_));
 sky130_fd_sc_hd__a21o_1 _08032_ (.A1(_07041_),
    .A2(_07073_),
    .B1(_07072_),
    .X(_00076_));
 sky130_fd_sc_hd__xor2_2 _08033_ (.A(_00075_),
    .B(_00076_),
    .X(_00077_));
 sky130_fd_sc_hd__and3_1 _08034_ (.A(_07039_),
    .B(_07075_),
    .C(_00077_),
    .X(_00078_));
 sky130_fd_sc_hd__a21oi_1 _08035_ (.A1(net165),
    .A2(_07075_),
    .B1(_00077_),
    .Y(_00079_));
 sky130_fd_sc_hd__or4_4 _08036_ (.A(_00041_),
    .B(_00042_),
    .C(_00078_),
    .D(_00079_),
    .X(_00080_));
 sky130_fd_sc_hd__buf_6 _08037_ (.A(_00080_),
    .X(_00081_));
 sky130_fd_sc_hd__o22ai_1 _08038_ (.A1(_00041_),
    .A2(_00042_),
    .B1(_00078_),
    .B2(_00079_),
    .Y(_00082_));
 sky130_fd_sc_hd__and3_1 _08039_ (.A(_00081_),
    .B(_07077_),
    .C(_00082_),
    .X(_00083_));
 sky130_fd_sc_hd__a21oi_1 _08040_ (.A1(_00081_),
    .A2(_00082_),
    .B1(_07077_),
    .Y(_00084_));
 sky130_fd_sc_hd__nor2_1 _08041_ (.A(_00083_),
    .B(_00084_),
    .Y(_00085_));
 sky130_fd_sc_hd__xnor2_1 _08042_ (.A(_00002_),
    .B(_00085_),
    .Y(_00086_));
 sky130_fd_sc_hd__nor2_1 _08043_ (.A(_07079_),
    .B(_07080_),
    .Y(_00087_));
 sky130_fd_sc_hd__a21boi_1 _08044_ (.A1(_07079_),
    .A2(_07080_),
    .B1_N(_07001_),
    .Y(_00088_));
 sky130_fd_sc_hd__or3_4 _08045_ (.A(_00086_),
    .B(_00087_),
    .C(_00088_),
    .X(_00089_));
 sky130_fd_sc_hd__o21ai_1 _08046_ (.A1(_00087_),
    .A2(_00088_),
    .B1(_00086_),
    .Y(_00090_));
 sky130_fd_sc_hd__and4_1 _08047_ (.A(_03521_),
    .B(_00377_),
    .C(_02982_),
    .D(_06875_),
    .X(_00091_));
 sky130_fd_sc_hd__a22o_1 _08048_ (.A1(_03521_),
    .A2(_02993_),
    .B1(_06875_),
    .B2(_00377_),
    .X(_00092_));
 sky130_fd_sc_hd__or2b_1 _08049_ (.A(_00091_),
    .B_N(_00092_),
    .X(_00093_));
 sky130_fd_sc_hd__clkbuf_4 _08050_ (.A(_05203_),
    .X(_00094_));
 sky130_fd_sc_hd__clkbuf_4 _08051_ (.A(_00094_),
    .X(_00095_));
 sky130_fd_sc_hd__nand2_1 _08052_ (.A(_00497_),
    .B(_00095_),
    .Y(_00096_));
 sky130_fd_sc_hd__xnor2_1 _08053_ (.A(_00093_),
    .B(_00096_),
    .Y(_00097_));
 sky130_fd_sc_hd__nor2_1 _08054_ (.A(_00000_),
    .B(_00097_),
    .Y(_00098_));
 sky130_fd_sc_hd__and2_1 _08055_ (.A(_00000_),
    .B(_00097_),
    .X(_00099_));
 sky130_fd_sc_hd__or2_2 _08056_ (.A(_00098_),
    .B(_00099_),
    .X(_00100_));
 sky130_fd_sc_hd__buf_2 _08057_ (.A(net38),
    .X(_00101_));
 sky130_fd_sc_hd__and4_1 _08058_ (.A(_00628_),
    .B(_00650_),
    .C(_00101_),
    .D(_06733_),
    .X(_00102_));
 sky130_fd_sc_hd__inv_2 _08059_ (.A(_00102_),
    .Y(_00103_));
 sky130_fd_sc_hd__a22o_1 _08060_ (.A1(_02105_),
    .A2(_00101_),
    .B1(_06733_),
    .B2(_00650_),
    .X(_00104_));
 sky130_fd_sc_hd__and4_1 _08061_ (.A(_05588_),
    .B(_06744_),
    .C(_00103_),
    .D(_00104_),
    .X(_00105_));
 sky130_fd_sc_hd__a22oi_1 _08062_ (.A1(_06472_),
    .A2(_06885_),
    .B1(_00103_),
    .B2(_00104_),
    .Y(_00106_));
 sky130_fd_sc_hd__nor2_1 _08063_ (.A(_00105_),
    .B(_00106_),
    .Y(_00107_));
 sky130_fd_sc_hd__nand2_1 _08064_ (.A(_00006_),
    .B(_00107_),
    .Y(_00108_));
 sky130_fd_sc_hd__or2_1 _08065_ (.A(_00006_),
    .B(_00107_),
    .X(_00109_));
 sky130_fd_sc_hd__nand2_1 _08066_ (.A(_00108_),
    .B(_00109_),
    .Y(_00110_));
 sky130_fd_sc_hd__and3_1 _08067_ (.A(_00009_),
    .B(_00010_),
    .C(_00011_),
    .X(_00111_));
 sky130_fd_sc_hd__clkbuf_4 _08068_ (.A(_07010_),
    .X(_00112_));
 sky130_fd_sc_hd__clkbuf_4 _08069_ (.A(_00112_),
    .X(_00113_));
 sky130_fd_sc_hd__clkbuf_4 _08070_ (.A(_00101_),
    .X(_00114_));
 sky130_fd_sc_hd__nand2_1 _08071_ (.A(_01383_),
    .B(_00114_),
    .Y(_00115_));
 sky130_fd_sc_hd__and3_1 _08072_ (.A(_01350_),
    .B(_00113_),
    .C(_00115_),
    .X(_00116_));
 sky130_fd_sc_hd__xor2_1 _08073_ (.A(_00111_),
    .B(_00116_),
    .X(_00117_));
 sky130_fd_sc_hd__o21ba_1 _08074_ (.A1(_00016_),
    .A2(_00018_),
    .B1_N(_00014_),
    .X(_00118_));
 sky130_fd_sc_hd__xnor2_1 _08075_ (.A(_00117_),
    .B(_00118_),
    .Y(_00119_));
 sky130_fd_sc_hd__and3_1 _08076_ (.A(_00021_),
    .B(_00022_),
    .C(_00023_),
    .X(_00120_));
 sky130_fd_sc_hd__clkbuf_4 _08077_ (.A(_06874_),
    .X(_00121_));
 sky130_fd_sc_hd__nand2_1 _08078_ (.A(_06461_),
    .B(_00121_),
    .Y(_00122_));
 sky130_fd_sc_hd__and3_1 _08079_ (.A(_05566_),
    .B(_06964_),
    .C(_00122_),
    .X(_00123_));
 sky130_fd_sc_hd__xor2_2 _08080_ (.A(_00120_),
    .B(_00123_),
    .X(_00124_));
 sky130_fd_sc_hd__o21ba_1 _08081_ (.A1(_00028_),
    .A2(_00030_),
    .B1_N(_00026_),
    .X(_00125_));
 sky130_fd_sc_hd__xnor2_2 _08082_ (.A(_00124_),
    .B(_00125_),
    .Y(_00126_));
 sky130_fd_sc_hd__xnor2_1 _08083_ (.A(_00119_),
    .B(_00126_),
    .Y(_00127_));
 sky130_fd_sc_hd__and2_1 _08084_ (.A(_00032_),
    .B(_00127_),
    .X(_00128_));
 sky130_fd_sc_hd__nor2_1 _08085_ (.A(_00032_),
    .B(_00127_),
    .Y(_00129_));
 sky130_fd_sc_hd__nor2_1 _08086_ (.A(_00128_),
    .B(_00129_),
    .Y(_00130_));
 sky130_fd_sc_hd__o21ai_1 _08087_ (.A1(_00032_),
    .A2(_00127_),
    .B1(_00110_),
    .Y(_00131_));
 sky130_fd_sc_hd__o22a_1 _08088_ (.A1(_00110_),
    .A2(_00130_),
    .B1(_00131_),
    .B2(_00128_),
    .X(_00132_));
 sky130_fd_sc_hd__a21bo_1 _08089_ (.A1(_00007_),
    .A2(_00036_),
    .B1_N(_00035_),
    .X(_00133_));
 sky130_fd_sc_hd__xnor2_2 _08090_ (.A(_00132_),
    .B(_00133_),
    .Y(_00134_));
 sky130_fd_sc_hd__nor2_1 _08091_ (.A(_00038_),
    .B(_00039_),
    .Y(_00135_));
 sky130_fd_sc_hd__a31o_1 _08092_ (.A1(_07003_),
    .A2(_07036_),
    .A3(_00040_),
    .B1(_00135_),
    .X(_00136_));
 sky130_fd_sc_hd__xnor2_1 _08093_ (.A(_00134_),
    .B(_00136_),
    .Y(_00137_));
 sky130_fd_sc_hd__buf_2 _08094_ (.A(_05478_),
    .X(_00138_));
 sky130_fd_sc_hd__and3_1 _08095_ (.A(_00138_),
    .B(_02007_),
    .C(_04928_),
    .X(_00139_));
 sky130_fd_sc_hd__a22o_1 _08096_ (.A1(_02018_),
    .A2(_04895_),
    .B1(_04928_),
    .B2(_05478_),
    .X(_00140_));
 sky130_fd_sc_hd__a21bo_1 _08097_ (.A1(_04917_),
    .A2(_00139_),
    .B1_N(_00140_),
    .X(_00141_));
 sky130_fd_sc_hd__clkbuf_4 _08098_ (.A(_05027_),
    .X(_00142_));
 sky130_fd_sc_hd__clkbuf_4 _08099_ (.A(_00142_),
    .X(_00143_));
 sky130_fd_sc_hd__clkbuf_4 _08100_ (.A(_00143_),
    .X(_00144_));
 sky130_fd_sc_hd__clkbuf_4 _08101_ (.A(_00144_),
    .X(_00145_));
 sky130_fd_sc_hd__nand2_1 _08102_ (.A(_02280_),
    .B(_00145_),
    .Y(_00146_));
 sky130_fd_sc_hd__xnor2_1 _08103_ (.A(_00141_),
    .B(_00146_),
    .Y(_00147_));
 sky130_fd_sc_hd__nor2_1 _08104_ (.A(_00045_),
    .B(_00147_),
    .Y(_00148_));
 sky130_fd_sc_hd__and2_1 _08105_ (.A(_00045_),
    .B(_00147_),
    .X(_00149_));
 sky130_fd_sc_hd__or2_1 _08106_ (.A(_00148_),
    .B(_00149_),
    .X(_00150_));
 sky130_fd_sc_hd__clkbuf_4 _08107_ (.A(_05181_),
    .X(_00151_));
 sky130_fd_sc_hd__nand2_1 _08108_ (.A(_05478_),
    .B(_00094_),
    .Y(_00152_));
 sky130_fd_sc_hd__and3_1 _08109_ (.A(_06417_),
    .B(_00151_),
    .C(_00152_),
    .X(_00153_));
 sky130_fd_sc_hd__xor2_1 _08110_ (.A(_00050_),
    .B(_00153_),
    .X(_00154_));
 sky130_fd_sc_hd__o21ba_1 _08111_ (.A1(_00055_),
    .A2(_00056_),
    .B1_N(_00053_),
    .X(_00155_));
 sky130_fd_sc_hd__xnor2_1 _08112_ (.A(_00154_),
    .B(_00155_),
    .Y(_00156_));
 sky130_fd_sc_hd__clkbuf_4 _08113_ (.A(_01361_),
    .X(_00157_));
 sky130_fd_sc_hd__clkbuf_4 _08114_ (.A(net7),
    .X(_00158_));
 sky130_fd_sc_hd__buf_4 _08115_ (.A(_01405_),
    .X(_00159_));
 sky130_fd_sc_hd__nand2_1 _08116_ (.A(_00159_),
    .B(_00142_),
    .Y(_00160_));
 sky130_fd_sc_hd__and3_1 _08117_ (.A(_00157_),
    .B(_00158_),
    .C(_00160_),
    .X(_00161_));
 sky130_fd_sc_hd__xor2_1 _08118_ (.A(_00061_),
    .B(_00161_),
    .X(_00162_));
 sky130_fd_sc_hd__o21ba_1 _08119_ (.A1(_00066_),
    .A2(_00067_),
    .B1_N(_00064_),
    .X(_00163_));
 sky130_fd_sc_hd__xnor2_1 _08120_ (.A(_00162_),
    .B(_00163_),
    .Y(_00164_));
 sky130_fd_sc_hd__xnor2_1 _08121_ (.A(_00156_),
    .B(_00164_),
    .Y(_00165_));
 sky130_fd_sc_hd__and2_1 _08122_ (.A(_00069_),
    .B(_00165_),
    .X(_00166_));
 sky130_fd_sc_hd__nor2_1 _08123_ (.A(_00069_),
    .B(_00165_),
    .Y(_00167_));
 sky130_fd_sc_hd__nor2_1 _08124_ (.A(_00166_),
    .B(_00167_),
    .Y(_00168_));
 sky130_fd_sc_hd__o21ai_1 _08125_ (.A1(_00069_),
    .A2(_00165_),
    .B1(_00150_),
    .Y(_00169_));
 sky130_fd_sc_hd__o22a_1 _08126_ (.A1(_00150_),
    .A2(_00168_),
    .B1(_00169_),
    .B2(_00166_),
    .X(_00170_));
 sky130_fd_sc_hd__a21bo_1 _08127_ (.A1(_00046_),
    .A2(_00073_),
    .B1_N(_00072_),
    .X(_00171_));
 sky130_fd_sc_hd__xnor2_2 _08128_ (.A(_00170_),
    .B(_00171_),
    .Y(_00172_));
 sky130_fd_sc_hd__nor2_1 _08129_ (.A(_00075_),
    .B(_00076_),
    .Y(_00173_));
 sky130_fd_sc_hd__a31o_2 _08130_ (.A1(_07039_),
    .A2(_07075_),
    .A3(_00077_),
    .B1(_00173_),
    .X(_00174_));
 sky130_fd_sc_hd__xnor2_2 _08131_ (.A(_00172_),
    .B(_00174_),
    .Y(_00175_));
 sky130_fd_sc_hd__xnor2_1 _08132_ (.A(_00137_),
    .B(_00175_),
    .Y(_00176_));
 sky130_fd_sc_hd__xor2_1 _08133_ (.A(_00081_),
    .B(_00176_),
    .X(_00177_));
 sky130_fd_sc_hd__xnor2_1 _08134_ (.A(_00100_),
    .B(_00177_),
    .Y(_00178_));
 sky130_fd_sc_hd__and2b_1 _08135_ (.A_N(_00084_),
    .B(_00002_),
    .X(_00179_));
 sky130_fd_sc_hd__nor3_2 _08136_ (.A(_00178_),
    .B(_00083_),
    .C(_00179_),
    .Y(_00180_));
 sky130_fd_sc_hd__o21ai_2 _08137_ (.A1(_00083_),
    .A2(_00179_),
    .B1(_00178_),
    .Y(_00181_));
 sky130_fd_sc_hd__and2b_1 _08138_ (.A_N(_00180_),
    .B(_00181_),
    .X(_00182_));
 sky130_fd_sc_hd__and3_1 _08139_ (.A(_00089_),
    .B(_00090_),
    .C(_00182_),
    .X(_00183_));
 sky130_fd_sc_hd__nand2_1 _08140_ (.A(_06985_),
    .B(_07082_),
    .Y(_00184_));
 sky130_fd_sc_hd__or2_1 _08141_ (.A(_06985_),
    .B(_07082_),
    .X(_00185_));
 sky130_fd_sc_hd__and2_1 _08142_ (.A(_00184_),
    .B(_00185_),
    .X(_00186_));
 sky130_fd_sc_hd__and2_1 _08143_ (.A(_06998_),
    .B(_06999_),
    .X(_00187_));
 sky130_fd_sc_hd__nor2_1 _08144_ (.A(_07000_),
    .B(_00187_),
    .Y(_00188_));
 sky130_fd_sc_hd__and3_1 _08145_ (.A(_00186_),
    .B(_00188_),
    .C(_00183_),
    .X(_00189_));
 sky130_fd_sc_hd__or3_4 _08146_ (.A(_06989_),
    .B(_06996_),
    .C(_06995_),
    .X(_00190_));
 sky130_fd_sc_hd__o21ai_1 _08147_ (.A1(_06996_),
    .A2(_06995_),
    .B1(_06989_),
    .Y(_00191_));
 sky130_fd_sc_hd__inv_2 _08148_ (.A(_05346_),
    .Y(_00192_));
 sky130_fd_sc_hd__nand2_1 _08149_ (.A(_05357_),
    .B(_00192_),
    .Y(_00193_));
 sky130_fd_sc_hd__xor2_2 _08150_ (.A(_05313_),
    .B(_00193_),
    .X(_00194_));
 sky130_fd_sc_hd__and3_1 _08151_ (.A(net150),
    .B(_06175_),
    .C(_06406_),
    .X(_00195_));
 sky130_fd_sc_hd__nor2_1 _08152_ (.A(_06990_),
    .B(_00195_),
    .Y(_00196_));
 sky130_fd_sc_hd__and2_1 _08153_ (.A(_06889_),
    .B(_06888_),
    .X(_00197_));
 sky130_fd_sc_hd__xnor2_2 _08154_ (.A(_06884_),
    .B(_00197_),
    .Y(_00198_));
 sky130_fd_sc_hd__nand2_1 _08155_ (.A(_00196_),
    .B(_00198_),
    .Y(_00199_));
 sky130_fd_sc_hd__nor2_1 _08156_ (.A(_00196_),
    .B(_00198_),
    .Y(_00200_));
 sky130_fd_sc_hd__a21o_1 _08157_ (.A1(_00194_),
    .A2(_00199_),
    .B1(_00200_),
    .X(_00201_));
 sky130_fd_sc_hd__a21oi_4 _08158_ (.A1(_00190_),
    .A2(_00191_),
    .B1(_00201_),
    .Y(_00202_));
 sky130_fd_sc_hd__nand3_1 _08159_ (.A(_06986_),
    .B(_06987_),
    .C(_06997_),
    .Y(_00203_));
 sky130_fd_sc_hd__and3_1 _08160_ (.A(_00202_),
    .B(_06998_),
    .C(_00203_),
    .X(_00204_));
 sky130_fd_sc_hd__a21oi_1 _08161_ (.A1(_06998_),
    .A2(_00203_),
    .B1(_00202_),
    .Y(_00205_));
 sky130_fd_sc_hd__or2_4 _08162_ (.A(_00204_),
    .B(_00205_),
    .X(_00206_));
 sky130_fd_sc_hd__nor2_1 _08163_ (.A(_04774_),
    .B(_04785_),
    .Y(_00207_));
 sky130_fd_sc_hd__nor2_2 _08164_ (.A(_04796_),
    .B(_00207_),
    .Y(_00208_));
 sky130_fd_sc_hd__nor2_1 _08165_ (.A(_06845_),
    .B(_06846_),
    .Y(_00209_));
 sky130_fd_sc_hd__or2_2 _08166_ (.A(_06847_),
    .B(_00209_),
    .X(_00210_));
 sky130_fd_sc_hd__or2b_1 _08167_ (.A(net167),
    .B_N(_06076_),
    .X(_00211_));
 sky130_fd_sc_hd__a31o_1 _08168_ (.A1(_02445_),
    .A2(_02883_),
    .A3(_03477_),
    .B1(net140),
    .X(_00212_));
 sky130_fd_sc_hd__a21oi_1 _08169_ (.A1(_06120_),
    .A2(_00212_),
    .B1(_06153_),
    .Y(_00213_));
 sky130_fd_sc_hd__xnor2_2 _08170_ (.A(_00211_),
    .B(_00213_),
    .Y(_00214_));
 sky130_fd_sc_hd__xnor2_1 _08171_ (.A(_00210_),
    .B(_00214_),
    .Y(_00215_));
 sky130_fd_sc_hd__xnor2_2 _08172_ (.A(_00208_),
    .B(_00215_),
    .Y(_00216_));
 sky130_fd_sc_hd__xnor2_2 _08173_ (.A(_06120_),
    .B(_00212_),
    .Y(_00217_));
 sky130_fd_sc_hd__nor2_1 _08174_ (.A(_03598_),
    .B(_06844_),
    .Y(_00218_));
 sky130_fd_sc_hd__or2_2 _08175_ (.A(_06845_),
    .B(_00218_),
    .X(_00219_));
 sky130_fd_sc_hd__nor2_1 _08176_ (.A(_03037_),
    .B(_04763_),
    .Y(_00220_));
 sky130_fd_sc_hd__nor2_1 _08177_ (.A(_04774_),
    .B(_00220_),
    .Y(_00221_));
 sky130_fd_sc_hd__o21ba_1 _08178_ (.A1(_00217_),
    .A2(_00219_),
    .B1_N(_00221_),
    .X(_00222_));
 sky130_fd_sc_hd__a21o_1 _08179_ (.A1(_00217_),
    .A2(_00219_),
    .B1(_00222_),
    .X(_00223_));
 sky130_fd_sc_hd__xnor2_2 _08180_ (.A(_00216_),
    .B(_00223_),
    .Y(_00224_));
 sky130_fd_sc_hd__a21bo_1 _08181_ (.A1(_03488_),
    .A2(_03609_),
    .B1_N(_03048_),
    .X(_00225_));
 sky130_fd_sc_hd__o21ai_4 _08182_ (.A1(_03488_),
    .A2(_03609_),
    .B1(_00225_),
    .Y(_00226_));
 sky130_fd_sc_hd__xor2_1 _08183_ (.A(_00217_),
    .B(_00219_),
    .X(_00227_));
 sky130_fd_sc_hd__xnor2_2 _08184_ (.A(_00221_),
    .B(_00227_),
    .Y(_00228_));
 sky130_fd_sc_hd__xnor2_4 _08185_ (.A(_00226_),
    .B(_00228_),
    .Y(_00229_));
 sky130_fd_sc_hd__and2b_1 _08186_ (.A_N(_00228_),
    .B(_00226_),
    .X(_00230_));
 sky130_fd_sc_hd__a31o_1 _08187_ (.A1(_02949_),
    .A2(_03631_),
    .A3(_00229_),
    .B1(_00230_),
    .X(_00231_));
 sky130_fd_sc_hd__and2b_1 _08188_ (.A_N(_00223_),
    .B(_00216_),
    .X(_00232_));
 sky130_fd_sc_hd__a21o_2 _08189_ (.A1(_00224_),
    .A2(_00231_),
    .B1(_00232_),
    .X(_00233_));
 sky130_fd_sc_hd__nand2_1 _08190_ (.A(_00210_),
    .B(_00214_),
    .Y(_00234_));
 sky130_fd_sc_hd__xor2_1 _08191_ (.A(_00196_),
    .B(_00198_),
    .X(_00235_));
 sky130_fd_sc_hd__xnor2_1 _08192_ (.A(_00194_),
    .B(_00235_),
    .Y(_00236_));
 sky130_fd_sc_hd__o21bai_1 _08193_ (.A1(_00210_),
    .A2(_00214_),
    .B1_N(_00208_),
    .Y(_00237_));
 sky130_fd_sc_hd__and3_1 _08194_ (.A(_00234_),
    .B(_00236_),
    .C(_00237_),
    .X(_00238_));
 sky130_fd_sc_hd__buf_2 _08195_ (.A(_00238_),
    .X(_00239_));
 sky130_fd_sc_hd__a21oi_1 _08196_ (.A1(_00234_),
    .A2(_00237_),
    .B1(_00236_),
    .Y(_00240_));
 sky130_fd_sc_hd__nor2_1 _08197_ (.A(_00239_),
    .B(_00240_),
    .Y(_00241_));
 sky130_fd_sc_hd__nand2_2 _08198_ (.A(_00233_),
    .B(_00241_),
    .Y(_00242_));
 sky130_fd_sc_hd__and3_1 _08199_ (.A(_00190_),
    .B(_00191_),
    .C(_00201_),
    .X(_00243_));
 sky130_fd_sc_hd__nor2_4 _08200_ (.A(_00202_),
    .B(_00243_),
    .Y(_00244_));
 sky130_fd_sc_hd__xnor2_2 _08201_ (.A(_00244_),
    .B(_00239_),
    .Y(_00245_));
 sky130_fd_sc_hd__a21oi_1 _08202_ (.A1(_00244_),
    .A2(_00239_),
    .B1(_00202_),
    .Y(_00246_));
 sky130_fd_sc_hd__and2_1 _08203_ (.A(_06998_),
    .B(_00203_),
    .X(_00247_));
 sky130_fd_sc_hd__inv_2 _08204_ (.A(_00247_),
    .Y(_00248_));
 sky130_fd_sc_hd__o32ai_4 _08205_ (.A1(_00206_),
    .A2(_00242_),
    .A3(_00245_),
    .B1(_00246_),
    .B2(_00248_),
    .Y(_00249_));
 sky130_fd_sc_hd__a21oi_1 _08206_ (.A1(_00089_),
    .A2(_00181_),
    .B1(_00180_),
    .Y(_00250_));
 sky130_fd_sc_hd__a221o_2 _08207_ (.A1(_07083_),
    .A2(_00183_),
    .B1(_00189_),
    .B2(_00249_),
    .C1(_00250_),
    .X(_00251_));
 sky130_fd_sc_hd__nor2_1 _08208_ (.A(_00081_),
    .B(_00176_),
    .Y(_00252_));
 sky130_fd_sc_hd__a21oi_1 _08209_ (.A1(_00081_),
    .A2(_00176_),
    .B1(_00100_),
    .Y(_00253_));
 sky130_fd_sc_hd__nor2_1 _08210_ (.A(_00137_),
    .B(_00175_),
    .Y(_00254_));
 sky130_fd_sc_hd__nand2_1 _08211_ (.A(_00119_),
    .B(_00126_),
    .Y(_00255_));
 sky130_fd_sc_hd__and2b_1 _08212_ (.A_N(_00118_),
    .B(_00117_),
    .X(_00256_));
 sky130_fd_sc_hd__clkbuf_4 _08213_ (.A(_00113_),
    .X(_00257_));
 sky130_fd_sc_hd__clkbuf_4 _08214_ (.A(_00114_),
    .X(_00258_));
 sky130_fd_sc_hd__and4_1 _08215_ (.A(_01383_),
    .B(_01350_),
    .C(_00257_),
    .D(_00258_),
    .X(_00259_));
 sky130_fd_sc_hd__a211o_1 _08216_ (.A1(_00111_),
    .A2(_00116_),
    .B1(_00256_),
    .C1(_00259_),
    .X(_00260_));
 sky130_fd_sc_hd__and2b_1 _08217_ (.A_N(_00125_),
    .B(_00124_),
    .X(_00261_));
 sky130_fd_sc_hd__clkbuf_4 _08218_ (.A(_06965_),
    .X(_00262_));
 sky130_fd_sc_hd__clkbuf_4 _08219_ (.A(_06966_),
    .X(_00263_));
 sky130_fd_sc_hd__and4_1 _08220_ (.A(_06472_),
    .B(_06483_),
    .C(_00262_),
    .D(_00263_),
    .X(_00264_));
 sky130_fd_sc_hd__a211o_2 _08221_ (.A1(_00120_),
    .A2(_00123_),
    .B1(_00261_),
    .C1(_00264_),
    .X(_00265_));
 sky130_fd_sc_hd__xnor2_2 _08222_ (.A(_00260_),
    .B(_00265_),
    .Y(_00266_));
 sky130_fd_sc_hd__xnor2_1 _08223_ (.A(_00255_),
    .B(_00266_),
    .Y(_00267_));
 sky130_fd_sc_hd__clkbuf_4 _08224_ (.A(_00101_),
    .X(_00268_));
 sky130_fd_sc_hd__and4_1 _08225_ (.A(_02116_),
    .B(_02149_),
    .C(_00112_),
    .D(_00268_),
    .X(_00269_));
 sky130_fd_sc_hd__a22o_1 _08226_ (.A1(_02116_),
    .A2(_00112_),
    .B1(_00268_),
    .B2(_02149_),
    .X(_00270_));
 sky130_fd_sc_hd__and2b_1 _08227_ (.A_N(_00269_),
    .B(_00270_),
    .X(_00271_));
 sky130_fd_sc_hd__nand2_1 _08228_ (.A(_06461_),
    .B(_00003_),
    .Y(_00272_));
 sky130_fd_sc_hd__xnor2_1 _08229_ (.A(_00271_),
    .B(_00272_),
    .Y(_00273_));
 sky130_fd_sc_hd__or2_1 _08230_ (.A(_00102_),
    .B(_00105_),
    .X(_00274_));
 sky130_fd_sc_hd__nand2_1 _08231_ (.A(_05566_),
    .B(_06775_),
    .Y(_00275_));
 sky130_fd_sc_hd__xnor2_1 _08232_ (.A(_00274_),
    .B(_00275_),
    .Y(_00276_));
 sky130_fd_sc_hd__and2_1 _08233_ (.A(_00273_),
    .B(_00276_),
    .X(_00277_));
 sky130_fd_sc_hd__nor2_1 _08234_ (.A(_00273_),
    .B(_00276_),
    .Y(_00278_));
 sky130_fd_sc_hd__or2_1 _08235_ (.A(_00277_),
    .B(_00278_),
    .X(_00279_));
 sky130_fd_sc_hd__nor2_1 _08236_ (.A(_00108_),
    .B(_00279_),
    .Y(_00280_));
 sky130_fd_sc_hd__and2_1 _08237_ (.A(_00108_),
    .B(_00279_),
    .X(_00281_));
 sky130_fd_sc_hd__or2_1 _08238_ (.A(_00280_),
    .B(_00281_),
    .X(_00282_));
 sky130_fd_sc_hd__xnor2_1 _08239_ (.A(_00267_),
    .B(_00282_),
    .Y(_00283_));
 sky130_fd_sc_hd__or2b_1 _08240_ (.A(_00128_),
    .B_N(_00131_),
    .X(_00284_));
 sky130_fd_sc_hd__and2_1 _08241_ (.A(_00283_),
    .B(_00284_),
    .X(_00285_));
 sky130_fd_sc_hd__nor2_1 _08242_ (.A(_00283_),
    .B(_00284_),
    .Y(_00286_));
 sky130_fd_sc_hd__nor2_1 _08243_ (.A(_00285_),
    .B(_00286_),
    .Y(_00287_));
 sky130_fd_sc_hd__and2b_1 _08244_ (.A_N(_00132_),
    .B(_00133_),
    .X(_00288_));
 sky130_fd_sc_hd__a21o_1 _08245_ (.A1(_00134_),
    .A2(_00136_),
    .B1(_00288_),
    .X(_00289_));
 sky130_fd_sc_hd__xnor2_2 _08246_ (.A(_00287_),
    .B(_00289_),
    .Y(_00290_));
 sky130_fd_sc_hd__nand2_1 _08247_ (.A(_00156_),
    .B(_00164_),
    .Y(_00291_));
 sky130_fd_sc_hd__and2b_1 _08248_ (.A_N(_00155_),
    .B(_00154_),
    .X(_00292_));
 sky130_fd_sc_hd__clkbuf_4 _08249_ (.A(_00095_),
    .X(_00293_));
 sky130_fd_sc_hd__clkbuf_4 _08250_ (.A(_00151_),
    .X(_00294_));
 sky130_fd_sc_hd__and4_1 _08251_ (.A(_06428_),
    .B(_06450_),
    .C(_00293_),
    .D(_00294_),
    .X(_00295_));
 sky130_fd_sc_hd__a211o_1 _08252_ (.A1(_00050_),
    .A2(_00153_),
    .B1(_00292_),
    .C1(_00295_),
    .X(_00296_));
 sky130_fd_sc_hd__and2b_1 _08253_ (.A_N(_00163_),
    .B(_00162_),
    .X(_00297_));
 sky130_fd_sc_hd__clkbuf_4 _08254_ (.A(_00158_),
    .X(_00298_));
 sky130_fd_sc_hd__and4_1 _08255_ (.A(_00157_),
    .B(_00159_),
    .C(_00144_),
    .D(_00298_),
    .X(_00299_));
 sky130_fd_sc_hd__a211o_1 _08256_ (.A1(_00061_),
    .A2(_00161_),
    .B1(_00297_),
    .C1(_00299_),
    .X(_00301_));
 sky130_fd_sc_hd__xnor2_2 _08257_ (.A(_00296_),
    .B(_00301_),
    .Y(_00302_));
 sky130_fd_sc_hd__xnor2_1 _08258_ (.A(_00291_),
    .B(_00302_),
    .Y(_00303_));
 sky130_fd_sc_hd__and4_1 _08259_ (.A(_06417_),
    .B(_00138_),
    .C(_04906_),
    .D(_04928_),
    .X(_00304_));
 sky130_fd_sc_hd__a22oi_1 _08260_ (.A1(_00138_),
    .A2(_04906_),
    .B1(_04928_),
    .B2(_06417_),
    .Y(_00305_));
 sky130_fd_sc_hd__and4bb_1 _08261_ (.A_N(_00304_),
    .B_N(_00305_),
    .C(_02018_),
    .D(_00143_),
    .X(_00306_));
 sky130_fd_sc_hd__o2bb2a_1 _08262_ (.A1_N(_03059_),
    .A2_N(_00144_),
    .B1(_00304_),
    .B2(_00305_),
    .X(_00307_));
 sky130_fd_sc_hd__a32o_1 _08263_ (.A1(_02040_),
    .A2(_00143_),
    .A3(_00140_),
    .B1(_00139_),
    .B2(_04917_),
    .X(_00308_));
 sky130_fd_sc_hd__and3_1 _08264_ (.A(_02040_),
    .B(_00298_),
    .C(_00308_),
    .X(_00309_));
 sky130_fd_sc_hd__clkbuf_4 _08265_ (.A(_00298_),
    .X(_00310_));
 sky130_fd_sc_hd__a21oi_1 _08266_ (.A1(_02280_),
    .A2(_00310_),
    .B1(_00308_),
    .Y(_00312_));
 sky130_fd_sc_hd__nor4_1 _08267_ (.A(_00306_),
    .B(_00307_),
    .C(_00309_),
    .D(_00312_),
    .Y(_00313_));
 sky130_fd_sc_hd__o22a_1 _08268_ (.A1(_00306_),
    .A2(_00307_),
    .B1(_00309_),
    .B2(_00312_),
    .X(_00314_));
 sky130_fd_sc_hd__nor2_1 _08269_ (.A(net145),
    .B(_00314_),
    .Y(_00315_));
 sky130_fd_sc_hd__nand2_1 _08270_ (.A(_00148_),
    .B(_00315_),
    .Y(_00316_));
 sky130_fd_sc_hd__or2_1 _08271_ (.A(_00148_),
    .B(_00315_),
    .X(_00317_));
 sky130_fd_sc_hd__nand2_1 _08272_ (.A(_00316_),
    .B(_00317_),
    .Y(_00318_));
 sky130_fd_sc_hd__xnor2_1 _08273_ (.A(_00303_),
    .B(_00318_),
    .Y(_00319_));
 sky130_fd_sc_hd__or2b_1 _08274_ (.A(_00166_),
    .B_N(_00169_),
    .X(_00320_));
 sky130_fd_sc_hd__and2_1 _08275_ (.A(_00319_),
    .B(_00320_),
    .X(_00321_));
 sky130_fd_sc_hd__nor2_1 _08276_ (.A(_00319_),
    .B(_00320_),
    .Y(_00323_));
 sky130_fd_sc_hd__nor2_2 _08277_ (.A(_00321_),
    .B(_00323_),
    .Y(_00324_));
 sky130_fd_sc_hd__and2b_1 _08278_ (.A_N(_00170_),
    .B(_00171_),
    .X(_00325_));
 sky130_fd_sc_hd__a21o_1 _08279_ (.A1(_00172_),
    .A2(_00174_),
    .B1(_00325_),
    .X(_00326_));
 sky130_fd_sc_hd__xnor2_4 _08280_ (.A(_00324_),
    .B(_00326_),
    .Y(_00327_));
 sky130_fd_sc_hd__xor2_2 _08281_ (.A(_00290_),
    .B(_00327_),
    .X(_00328_));
 sky130_fd_sc_hd__xor2_1 _08282_ (.A(_00254_),
    .B(_00328_),
    .X(_00329_));
 sky130_fd_sc_hd__and4_1 _08283_ (.A(_00377_),
    .B(_02982_),
    .C(_06873_),
    .D(_06874_),
    .X(_00330_));
 sky130_fd_sc_hd__a22o_1 _08284_ (.A1(_00377_),
    .A2(_06873_),
    .B1(_06875_),
    .B2(_02993_),
    .X(_00331_));
 sky130_fd_sc_hd__or2b_1 _08285_ (.A(_00330_),
    .B_N(_00331_),
    .X(_00332_));
 sky130_fd_sc_hd__nand2_1 _08286_ (.A(_03532_),
    .B(_00094_),
    .Y(_00334_));
 sky130_fd_sc_hd__xnor2_1 _08287_ (.A(_00332_),
    .B(_00334_),
    .Y(_00335_));
 sky130_fd_sc_hd__a31o_1 _08288_ (.A1(_00497_),
    .A2(_00094_),
    .A3(_00092_),
    .B1(_00091_),
    .X(_00336_));
 sky130_fd_sc_hd__nand2_1 _08289_ (.A(_00497_),
    .B(_00151_),
    .Y(_00337_));
 sky130_fd_sc_hd__xnor2_1 _08290_ (.A(_00336_),
    .B(_00337_),
    .Y(_00338_));
 sky130_fd_sc_hd__xnor2_1 _08291_ (.A(_00335_),
    .B(_00338_),
    .Y(_00339_));
 sky130_fd_sc_hd__nand2_2 _08292_ (.A(_00098_),
    .B(_00339_),
    .Y(_00340_));
 sky130_fd_sc_hd__or2_1 _08293_ (.A(_00098_),
    .B(_00339_),
    .X(_00341_));
 sky130_fd_sc_hd__nand2_1 _08294_ (.A(_00340_),
    .B(_00341_),
    .Y(_00342_));
 sky130_fd_sc_hd__xnor2_1 _08295_ (.A(_00329_),
    .B(_00342_),
    .Y(_00343_));
 sky130_fd_sc_hd__o21a_1 _08296_ (.A1(_00252_),
    .A2(_00253_),
    .B1(_00343_),
    .X(_00345_));
 sky130_fd_sc_hd__nor3_1 _08297_ (.A(_00252_),
    .B(_00253_),
    .C(_00343_),
    .Y(_00346_));
 sky130_fd_sc_hd__nor2_1 _08298_ (.A(_00345_),
    .B(_00346_),
    .Y(_00347_));
 sky130_fd_sc_hd__xnor2_4 _08299_ (.A(_00251_),
    .B(_00347_),
    .Y(_00348_));
 sky130_fd_sc_hd__xor2_2 _08300_ (.A(_04334_),
    .B(_00348_),
    .X(_00349_));
 sky130_fd_sc_hd__xnor2_4 _08301_ (.A(_04004_),
    .B(_00349_),
    .Y(_00350_));
 sky130_fd_sc_hd__or2_1 _08302_ (.A(_03751_),
    .B(_03828_),
    .X(_00351_));
 sky130_fd_sc_hd__and2_2 _08303_ (.A(_03839_),
    .B(_00351_),
    .X(_00352_));
 sky130_fd_sc_hd__or2_1 _08304_ (.A(_04070_),
    .B(_04147_),
    .X(_00353_));
 sky130_fd_sc_hd__nand2_2 _08305_ (.A(_04158_),
    .B(_00353_),
    .Y(_00354_));
 sky130_fd_sc_hd__xnor2_1 _08306_ (.A(_06985_),
    .B(_07082_),
    .Y(_00356_));
 sky130_fd_sc_hd__nand2_1 _08307_ (.A(_00089_),
    .B(_00090_),
    .Y(_00357_));
 sky130_fd_sc_hd__or2_1 _08308_ (.A(_00356_),
    .B(_00357_),
    .X(_00358_));
 sky130_fd_sc_hd__inv_2 _08309_ (.A(_00240_),
    .Y(_00359_));
 sky130_fd_sc_hd__o211ai_4 _08310_ (.A1(_00233_),
    .A2(_00239_),
    .B1(_00359_),
    .C1(_00244_),
    .Y(_00360_));
 sky130_fd_sc_hd__xnor2_2 _08311_ (.A(_06998_),
    .B(_06999_),
    .Y(_00361_));
 sky130_fd_sc_hd__or3_4 _08312_ (.A(_00204_),
    .B(_00205_),
    .C(_00361_),
    .X(_00362_));
 sky130_fd_sc_hd__a21boi_1 _08313_ (.A1(_00202_),
    .A2(_00203_),
    .B1_N(_06998_),
    .Y(_00363_));
 sky130_fd_sc_hd__or4_4 _08314_ (.A(_00356_),
    .B(_06999_),
    .C(_00357_),
    .D(_00363_),
    .X(_00364_));
 sky130_fd_sc_hd__a21bo_1 _08315_ (.A1(_00089_),
    .A2(_00184_),
    .B1_N(_00090_),
    .X(_00365_));
 sky130_fd_sc_hd__o311a_4 _08316_ (.A1(_00358_),
    .A2(_00360_),
    .A3(_00362_),
    .B1(_00364_),
    .C1(_00365_),
    .X(_00367_));
 sky130_fd_sc_hd__xor2_2 _08317_ (.A(net182),
    .B(_00367_),
    .X(_00368_));
 sky130_fd_sc_hd__nor2_1 _08318_ (.A(_00354_),
    .B(_00368_),
    .Y(_00369_));
 sky130_fd_sc_hd__nand2_1 _08319_ (.A(_00354_),
    .B(_00368_),
    .Y(_00370_));
 sky130_fd_sc_hd__o21ai_2 _08320_ (.A1(_00352_),
    .A2(_00369_),
    .B1(_00370_),
    .Y(_00371_));
 sky130_fd_sc_hd__xnor2_4 _08321_ (.A(_00350_),
    .B(_00371_),
    .Y(_00372_));
 sky130_fd_sc_hd__clkbuf_4 _08322_ (.A(_04015_),
    .X(_00373_));
 sky130_fd_sc_hd__clkbuf_4 _08323_ (.A(_00373_),
    .X(_00374_));
 sky130_fd_sc_hd__clkbuf_4 _08324_ (.A(_00374_),
    .X(_00375_));
 sky130_fd_sc_hd__buf_4 _08325_ (.A(_00375_),
    .X(_00376_));
 sky130_fd_sc_hd__clkbuf_4 _08326_ (.A(_04059_),
    .X(_00378_));
 sky130_fd_sc_hd__clkbuf_4 _08327_ (.A(_00378_),
    .X(_00379_));
 sky130_fd_sc_hd__clkbuf_8 _08328_ (.A(_00379_),
    .X(_00380_));
 sky130_fd_sc_hd__clkbuf_8 _08329_ (.A(_00380_),
    .X(_00381_));
 sky130_fd_sc_hd__a22oi_1 _08330_ (.A1(_00464_),
    .A2(_00376_),
    .B1(_00381_),
    .B2(_02051_),
    .Y(_00382_));
 sky130_fd_sc_hd__or2_1 _08331_ (.A(_04070_),
    .B(_00382_),
    .X(_00383_));
 sky130_fd_sc_hd__inv_2 _08332_ (.A(_00383_),
    .Y(_00384_));
 sky130_fd_sc_hd__a31o_1 _08333_ (.A1(_00186_),
    .A2(_00249_),
    .A3(_00188_),
    .B1(_07083_),
    .X(_00385_));
 sky130_fd_sc_hd__xnor2_2 _08334_ (.A(_00385_),
    .B(_00357_),
    .Y(_00386_));
 sky130_fd_sc_hd__and2_1 _08335_ (.A(_00384_),
    .B(_00386_),
    .X(_00387_));
 sky130_fd_sc_hd__clkbuf_4 _08336_ (.A(_03707_),
    .X(_00389_));
 sky130_fd_sc_hd__buf_4 _08337_ (.A(_00389_),
    .X(_00390_));
 sky130_fd_sc_hd__buf_6 _08338_ (.A(_00390_),
    .X(_00391_));
 sky130_fd_sc_hd__buf_4 _08339_ (.A(_03740_),
    .X(_00392_));
 sky130_fd_sc_hd__buf_4 _08340_ (.A(_00392_),
    .X(_00393_));
 sky130_fd_sc_hd__a22oi_1 _08341_ (.A1(_02138_),
    .A2(_00391_),
    .B1(_00393_),
    .B2(_00344_),
    .Y(_00394_));
 sky130_fd_sc_hd__nor2_2 _08342_ (.A(_03751_),
    .B(_00394_),
    .Y(_00395_));
 sky130_fd_sc_hd__o21a_1 _08343_ (.A1(_00384_),
    .A2(_00386_),
    .B1(_00395_),
    .X(_00396_));
 sky130_fd_sc_hd__xnor2_1 _08344_ (.A(_00354_),
    .B(_00368_),
    .Y(_00397_));
 sky130_fd_sc_hd__xnor2_1 _08345_ (.A(_00352_),
    .B(_00397_),
    .Y(_00398_));
 sky130_fd_sc_hd__or3_1 _08346_ (.A(_00387_),
    .B(_00396_),
    .C(_00398_),
    .X(_00400_));
 sky130_fd_sc_hd__and2_1 _08347_ (.A(_00344_),
    .B(_00391_),
    .X(_00401_));
 sky130_fd_sc_hd__o22a_1 _08348_ (.A1(_06999_),
    .A2(_00363_),
    .B1(_00360_),
    .B2(_00362_),
    .X(_00402_));
 sky130_fd_sc_hd__xnor2_1 _08349_ (.A(_00186_),
    .B(_00402_),
    .Y(_00403_));
 sky130_fd_sc_hd__and3_1 _08350_ (.A(_00464_),
    .B(_00381_),
    .C(_00403_),
    .X(_00404_));
 sky130_fd_sc_hd__a21o_1 _08351_ (.A1(_00464_),
    .A2(_00381_),
    .B1(_00403_),
    .X(_00405_));
 sky130_fd_sc_hd__o21a_1 _08352_ (.A1(_00401_),
    .A2(_00404_),
    .B1(_00405_),
    .X(_00406_));
 sky130_fd_sc_hd__xnor2_1 _08353_ (.A(_00384_),
    .B(_00386_),
    .Y(_00407_));
 sky130_fd_sc_hd__xnor2_1 _08354_ (.A(_00395_),
    .B(_00407_),
    .Y(_00408_));
 sky130_fd_sc_hd__o21a_1 _08355_ (.A1(_00387_),
    .A2(_00396_),
    .B1(_00398_),
    .X(_00409_));
 sky130_fd_sc_hd__a31o_2 _08356_ (.A1(_00400_),
    .A2(_00406_),
    .A3(_00408_),
    .B1(_00409_),
    .X(_00411_));
 sky130_fd_sc_hd__xor2_2 _08357_ (.A(_00372_),
    .B(_00411_),
    .X(net75));
 sky130_fd_sc_hd__nand2_1 _08358_ (.A(_04334_),
    .B(_00348_),
    .Y(_00412_));
 sky130_fd_sc_hd__buf_2 _08359_ (.A(net13),
    .X(_00413_));
 sky130_fd_sc_hd__clkbuf_4 _08360_ (.A(_00413_),
    .X(_00414_));
 sky130_fd_sc_hd__clkbuf_4 _08361_ (.A(_00414_),
    .X(_00415_));
 sky130_fd_sc_hd__buf_4 _08362_ (.A(_00415_),
    .X(_00416_));
 sky130_fd_sc_hd__nand2_2 _08363_ (.A(_00333_),
    .B(_00416_),
    .Y(_00417_));
 sky130_fd_sc_hd__or2b_1 _08364_ (.A(_03949_),
    .B_N(_03927_),
    .X(_00418_));
 sky130_fd_sc_hd__nand2_1 _08365_ (.A(_03916_),
    .B(_03960_),
    .Y(_00419_));
 sky130_fd_sc_hd__a31o_1 _08366_ (.A1(_02127_),
    .A2(_03894_),
    .A3(_03872_),
    .B1(_03861_),
    .X(_00421_));
 sky130_fd_sc_hd__and4_1 _08367_ (.A(_03850_),
    .B(_04510_),
    .C(net9),
    .D(net10),
    .X(_00422_));
 sky130_fd_sc_hd__clkbuf_4 _08368_ (.A(net9),
    .X(_00423_));
 sky130_fd_sc_hd__a22oi_1 _08369_ (.A1(_03850_),
    .A2(_00423_),
    .B1(net10),
    .B2(_01306_),
    .Y(_00424_));
 sky130_fd_sc_hd__and4bb_1 _08370_ (.A_N(_00422_),
    .B_N(_00424_),
    .C(_00672_),
    .D(net11),
    .X(_00425_));
 sky130_fd_sc_hd__o2bb2a_1 _08371_ (.A1_N(_01744_),
    .A2_N(net11),
    .B1(_00422_),
    .B2(_00424_),
    .X(_00426_));
 sky130_fd_sc_hd__nor2_1 _08372_ (.A(_00425_),
    .B(_00426_),
    .Y(_00427_));
 sky130_fd_sc_hd__xnor2_1 _08373_ (.A(_00421_),
    .B(_00427_),
    .Y(_00428_));
 sky130_fd_sc_hd__a21o_1 _08374_ (.A1(_00418_),
    .A2(_00419_),
    .B1(_00428_),
    .X(_00429_));
 sky130_fd_sc_hd__nand3_1 _08375_ (.A(_00418_),
    .B(_00419_),
    .C(_00428_),
    .Y(_00430_));
 sky130_fd_sc_hd__and3_1 _08376_ (.A(_03982_),
    .B(_00429_),
    .C(_00430_),
    .X(_00432_));
 sky130_fd_sc_hd__a21oi_1 _08377_ (.A1(_00429_),
    .A2(_00430_),
    .B1(_03982_),
    .Y(_00433_));
 sky130_fd_sc_hd__nor2_1 _08378_ (.A(_00432_),
    .B(_00433_),
    .Y(_00434_));
 sky130_fd_sc_hd__and2_1 _08379_ (.A(_02335_),
    .B(_00389_),
    .X(_00435_));
 sky130_fd_sc_hd__nand2_1 _08380_ (.A(_00434_),
    .B(_00435_),
    .Y(_00436_));
 sky130_fd_sc_hd__or2_1 _08381_ (.A(_00434_),
    .B(_00435_),
    .X(_00437_));
 sky130_fd_sc_hd__and2_1 _08382_ (.A(_00436_),
    .B(_00437_),
    .X(_00438_));
 sky130_fd_sc_hd__xor2_4 _08383_ (.A(_00417_),
    .B(_00438_),
    .X(_00439_));
 sky130_fd_sc_hd__nand2_1 _08384_ (.A(_02467_),
    .B(_00381_),
    .Y(_00440_));
 sky130_fd_sc_hd__or2b_1 _08385_ (.A(_04279_),
    .B_N(_04257_),
    .X(_00441_));
 sky130_fd_sc_hd__nand2_1 _08386_ (.A(_04246_),
    .B(_04290_),
    .Y(_00443_));
 sky130_fd_sc_hd__a31o_1 _08387_ (.A1(_04081_),
    .A2(_00373_),
    .A3(_04213_),
    .B1(_04202_),
    .X(_00444_));
 sky130_fd_sc_hd__and4_1 _08388_ (.A(_00978_),
    .B(_00880_),
    .C(_04180_),
    .D(net43),
    .X(_00445_));
 sky130_fd_sc_hd__a22o_1 _08389_ (.A1(_00880_),
    .A2(_04180_),
    .B1(_04191_),
    .B2(_04169_),
    .X(_00446_));
 sky130_fd_sc_hd__and2b_1 _08390_ (.A_N(_00445_),
    .B(_00446_),
    .X(_00447_));
 sky130_fd_sc_hd__nand2_1 _08391_ (.A(_04268_),
    .B(_04026_),
    .Y(_00448_));
 sky130_fd_sc_hd__xnor2_1 _08392_ (.A(_00447_),
    .B(_00448_),
    .Y(_00449_));
 sky130_fd_sc_hd__xnor2_1 _08393_ (.A(_00444_),
    .B(_00449_),
    .Y(_00450_));
 sky130_fd_sc_hd__a21o_1 _08394_ (.A1(_00441_),
    .A2(_00443_),
    .B1(_00450_),
    .X(_00451_));
 sky130_fd_sc_hd__nand3_1 _08395_ (.A(_00441_),
    .B(_00443_),
    .C(_00450_),
    .Y(_00452_));
 sky130_fd_sc_hd__and3_1 _08396_ (.A(_04312_),
    .B(_00451_),
    .C(_00452_),
    .X(_00454_));
 sky130_fd_sc_hd__a21oi_1 _08397_ (.A1(_00451_),
    .A2(_00452_),
    .B1(_04312_),
    .Y(_00455_));
 sky130_fd_sc_hd__nor2_1 _08398_ (.A(_00454_),
    .B(_00455_),
    .Y(_00456_));
 sky130_fd_sc_hd__clkbuf_4 _08399_ (.A(net45),
    .X(_00457_));
 sky130_fd_sc_hd__clkbuf_4 _08400_ (.A(_00457_),
    .X(_00458_));
 sky130_fd_sc_hd__buf_4 _08401_ (.A(_00458_),
    .X(_00459_));
 sky130_fd_sc_hd__buf_4 _08402_ (.A(_00459_),
    .X(_00460_));
 sky130_fd_sc_hd__nand2_1 _08403_ (.A(_00453_),
    .B(_00460_),
    .Y(_00461_));
 sky130_fd_sc_hd__xnor2_1 _08404_ (.A(_00456_),
    .B(_00461_),
    .Y(_00462_));
 sky130_fd_sc_hd__xnor2_1 _08405_ (.A(_00440_),
    .B(_00462_),
    .Y(_00463_));
 sky130_fd_sc_hd__nor2_1 _08406_ (.A(_00254_),
    .B(_00328_),
    .Y(_00465_));
 sky130_fd_sc_hd__nor2_1 _08407_ (.A(_00290_),
    .B(_00327_),
    .Y(_00466_));
 sky130_fd_sc_hd__nand2_1 _08408_ (.A(_00283_),
    .B(_00284_),
    .Y(_00467_));
 sky130_fd_sc_hd__a21o_1 _08409_ (.A1(_00288_),
    .A2(_00467_),
    .B1(_00286_),
    .X(_00468_));
 sky130_fd_sc_hd__a31o_1 _08410_ (.A1(_00134_),
    .A2(_00136_),
    .A3(_00287_),
    .B1(_00468_),
    .X(_00469_));
 sky130_fd_sc_hd__a31o_1 _08411_ (.A1(_06494_),
    .A2(_07004_),
    .A3(_00274_),
    .B1(_00277_),
    .X(_00470_));
 sky130_fd_sc_hd__a22o_1 _08412_ (.A1(_02149_),
    .A2(_00112_),
    .B1(_00268_),
    .B2(_05588_),
    .X(_00471_));
 sky130_fd_sc_hd__and4_1 _08413_ (.A(_02149_),
    .B(_05577_),
    .C(_07010_),
    .D(_00101_),
    .X(_00472_));
 sky130_fd_sc_hd__inv_2 _08414_ (.A(_00472_),
    .Y(_00473_));
 sky130_fd_sc_hd__and2_1 _08415_ (.A(_00471_),
    .B(_00473_),
    .X(_00474_));
 sky130_fd_sc_hd__nand2_1 _08416_ (.A(_06483_),
    .B(_00003_),
    .Y(_00476_));
 sky130_fd_sc_hd__xor2_1 _08417_ (.A(_00474_),
    .B(_00476_),
    .X(_00477_));
 sky130_fd_sc_hd__a31o_1 _08418_ (.A1(_06472_),
    .A2(_00003_),
    .A3(_00270_),
    .B1(_00269_),
    .X(_00478_));
 sky130_fd_sc_hd__and2b_1 _08419_ (.A_N(_00477_),
    .B(_00478_),
    .X(_00479_));
 sky130_fd_sc_hd__and2b_1 _08420_ (.A_N(_00478_),
    .B(_00477_),
    .X(_00480_));
 sky130_fd_sc_hd__or2_1 _08421_ (.A(_00479_),
    .B(_00480_),
    .X(_00481_));
 sky130_fd_sc_hd__xnor2_1 _08422_ (.A(_00470_),
    .B(_00481_),
    .Y(_00482_));
 sky130_fd_sc_hd__xnor2_1 _08423_ (.A(_00280_),
    .B(_00482_),
    .Y(_00483_));
 sky130_fd_sc_hd__and3b_1 _08424_ (.A_N(_00483_),
    .B(_00265_),
    .C(_00260_),
    .X(_00484_));
 sky130_fd_sc_hd__a21boi_1 _08425_ (.A1(_00260_),
    .A2(_00265_),
    .B1_N(_00483_),
    .Y(_00485_));
 sky130_fd_sc_hd__or2_1 _08426_ (.A(_00484_),
    .B(_00485_),
    .X(_00487_));
 sky130_fd_sc_hd__o21a_1 _08427_ (.A1(_00255_),
    .A2(_00266_),
    .B1(_00282_),
    .X(_00488_));
 sky130_fd_sc_hd__a21o_1 _08428_ (.A1(_00255_),
    .A2(_00266_),
    .B1(_00488_),
    .X(_00489_));
 sky130_fd_sc_hd__nor2_1 _08429_ (.A(_00487_),
    .B(_00489_),
    .Y(_00490_));
 sky130_fd_sc_hd__and2_1 _08430_ (.A(_00487_),
    .B(_00489_),
    .X(_00491_));
 sky130_fd_sc_hd__nor2_2 _08431_ (.A(_00490_),
    .B(_00491_),
    .Y(_00492_));
 sky130_fd_sc_hd__xnor2_2 _08432_ (.A(_00469_),
    .B(_00492_),
    .Y(_00493_));
 sky130_fd_sc_hd__nand2_1 _08433_ (.A(_00319_),
    .B(_00320_),
    .Y(_00494_));
 sky130_fd_sc_hd__a21o_1 _08434_ (.A1(_00325_),
    .A2(_00494_),
    .B1(_00323_),
    .X(_00495_));
 sky130_fd_sc_hd__a31o_2 _08435_ (.A1(_00172_),
    .A2(_00174_),
    .A3(_00324_),
    .B1(_00495_),
    .X(_00496_));
 sky130_fd_sc_hd__nand2_1 _08436_ (.A(_05478_),
    .B(_00142_),
    .Y(_00498_));
 sky130_fd_sc_hd__a21boi_1 _08437_ (.A1(_05456_),
    .A2(_04895_),
    .B1_N(_00498_),
    .Y(_00499_));
 sky130_fd_sc_hd__and4_1 _08438_ (.A(_05456_),
    .B(_05478_),
    .C(_00142_),
    .D(_04862_),
    .X(_00500_));
 sky130_fd_sc_hd__nor2_1 _08439_ (.A(_00499_),
    .B(_00500_),
    .Y(_00501_));
 sky130_fd_sc_hd__and3_1 _08440_ (.A(_02018_),
    .B(_00158_),
    .C(_00501_),
    .X(_00502_));
 sky130_fd_sc_hd__a21oi_1 _08441_ (.A1(_03059_),
    .A2(_00158_),
    .B1(_00501_),
    .Y(_00503_));
 sky130_fd_sc_hd__nor2_1 _08442_ (.A(_00502_),
    .B(_00503_),
    .Y(_00504_));
 sky130_fd_sc_hd__o21a_1 _08443_ (.A1(_00304_),
    .A2(_00306_),
    .B1(_00504_),
    .X(_00505_));
 sky130_fd_sc_hd__nor3_1 _08444_ (.A(_00304_),
    .B(_00306_),
    .C(_00504_),
    .Y(_00506_));
 sky130_fd_sc_hd__nor2_1 _08445_ (.A(_00505_),
    .B(_00506_),
    .Y(_00507_));
 sky130_fd_sc_hd__o21a_1 _08446_ (.A1(_00309_),
    .A2(net145),
    .B1(_00507_),
    .X(_00509_));
 sky130_fd_sc_hd__nor3_1 _08447_ (.A(_00309_),
    .B(_00313_),
    .C(_00507_),
    .Y(_00510_));
 sky130_fd_sc_hd__nor2_1 _08448_ (.A(_00509_),
    .B(_00510_),
    .Y(_00511_));
 sky130_fd_sc_hd__xnor2_1 _08449_ (.A(_00316_),
    .B(_00511_),
    .Y(_00512_));
 sky130_fd_sc_hd__and3_2 _08450_ (.A(_00296_),
    .B(_00301_),
    .C(_00512_),
    .X(_00513_));
 sky130_fd_sc_hd__and2_1 _08451_ (.A(_00296_),
    .B(_00301_),
    .X(_00514_));
 sky130_fd_sc_hd__nor2_1 _08452_ (.A(_00514_),
    .B(_00512_),
    .Y(_00515_));
 sky130_fd_sc_hd__or2_1 _08453_ (.A(_00513_),
    .B(_00515_),
    .X(_00516_));
 sky130_fd_sc_hd__o21a_1 _08454_ (.A1(_00291_),
    .A2(_00302_),
    .B1(_00318_),
    .X(_00517_));
 sky130_fd_sc_hd__a21o_1 _08455_ (.A1(_00291_),
    .A2(_00302_),
    .B1(_00517_),
    .X(_00518_));
 sky130_fd_sc_hd__nor2_1 _08456_ (.A(_00516_),
    .B(_00518_),
    .Y(_00520_));
 sky130_fd_sc_hd__and2_1 _08457_ (.A(_00516_),
    .B(_00518_),
    .X(_00521_));
 sky130_fd_sc_hd__nor2_2 _08458_ (.A(_00520_),
    .B(_00521_),
    .Y(_00522_));
 sky130_fd_sc_hd__xnor2_4 _08459_ (.A(_00496_),
    .B(_00522_),
    .Y(_00523_));
 sky130_fd_sc_hd__xor2_2 _08460_ (.A(_00493_),
    .B(_00523_),
    .X(_00524_));
 sky130_fd_sc_hd__xor2_1 _08461_ (.A(_00466_),
    .B(_00524_),
    .X(_00525_));
 sky130_fd_sc_hd__buf_4 _08462_ (.A(_07040_),
    .X(_00526_));
 sky130_fd_sc_hd__nand2_1 _08463_ (.A(_00519_),
    .B(_00526_),
    .Y(_00527_));
 sky130_fd_sc_hd__and3_1 _08464_ (.A(_00508_),
    .B(_00294_),
    .C(_00336_),
    .X(_00528_));
 sky130_fd_sc_hd__and2b_1 _08465_ (.A_N(_00335_),
    .B(_00338_),
    .X(_00529_));
 sky130_fd_sc_hd__a31o_1 _08466_ (.A1(_03543_),
    .A2(_00095_),
    .A3(_00331_),
    .B1(_00330_),
    .X(_00531_));
 sky130_fd_sc_hd__and4_1 _08467_ (.A(_02993_),
    .B(_06873_),
    .C(_06875_),
    .D(_05203_),
    .X(_00532_));
 sky130_fd_sc_hd__a22o_1 _08468_ (.A1(_02993_),
    .A2(_06873_),
    .B1(_06875_),
    .B2(_05203_),
    .X(_00533_));
 sky130_fd_sc_hd__and2b_1 _08469_ (.A_N(_00532_),
    .B(_00533_),
    .X(_00534_));
 sky130_fd_sc_hd__nand2_1 _08470_ (.A(_03532_),
    .B(_00151_),
    .Y(_00535_));
 sky130_fd_sc_hd__xnor2_1 _08471_ (.A(_00534_),
    .B(_00535_),
    .Y(_00536_));
 sky130_fd_sc_hd__xor2_1 _08472_ (.A(_00531_),
    .B(_00536_),
    .X(_00537_));
 sky130_fd_sc_hd__o21a_1 _08473_ (.A1(_00528_),
    .A2(_00529_),
    .B1(_00537_),
    .X(_00538_));
 sky130_fd_sc_hd__nor3_1 _08474_ (.A(_00528_),
    .B(_00529_),
    .C(_00537_),
    .Y(_00539_));
 sky130_fd_sc_hd__nor2_1 _08475_ (.A(_00538_),
    .B(_00539_),
    .Y(_00540_));
 sky130_fd_sc_hd__xnor2_2 _08476_ (.A(_00340_),
    .B(_00540_),
    .Y(_00542_));
 sky130_fd_sc_hd__buf_4 _08477_ (.A(_07004_),
    .X(_00543_));
 sky130_fd_sc_hd__buf_4 _08478_ (.A(_00543_),
    .X(_00544_));
 sky130_fd_sc_hd__nand2_1 _08479_ (.A(_00399_),
    .B(_00544_),
    .Y(_00545_));
 sky130_fd_sc_hd__xnor2_1 _08480_ (.A(_00542_),
    .B(_00545_),
    .Y(_00546_));
 sky130_fd_sc_hd__xnor2_2 _08481_ (.A(_00527_),
    .B(_00546_),
    .Y(_00547_));
 sky130_fd_sc_hd__xnor2_1 _08482_ (.A(_00525_),
    .B(_00547_),
    .Y(_00548_));
 sky130_fd_sc_hd__a21boi_1 _08483_ (.A1(_00254_),
    .A2(_00328_),
    .B1_N(_00342_),
    .Y(_00549_));
 sky130_fd_sc_hd__nor3_1 _08484_ (.A(_00465_),
    .B(_00548_),
    .C(_00549_),
    .Y(_00550_));
 sky130_fd_sc_hd__o21a_1 _08485_ (.A1(_00465_),
    .A2(_00549_),
    .B1(_00548_),
    .X(_00551_));
 sky130_fd_sc_hd__or2_1 _08486_ (.A(_00550_),
    .B(_00551_),
    .X(_00553_));
 sky130_fd_sc_hd__nand2_1 _08487_ (.A(net182),
    .B(_00347_),
    .Y(_00554_));
 sky130_fd_sc_hd__o21ai_1 _08488_ (.A1(_00252_),
    .A2(_00253_),
    .B1(_00343_),
    .Y(_00555_));
 sky130_fd_sc_hd__a21o_1 _08489_ (.A1(_00181_),
    .A2(_00555_),
    .B1(_00346_),
    .X(_00556_));
 sky130_fd_sc_hd__o21ai_4 _08490_ (.A1(_00367_),
    .A2(_00554_),
    .B1(_00556_),
    .Y(_00557_));
 sky130_fd_sc_hd__xnor2_2 _08491_ (.A(_00553_),
    .B(_00557_),
    .Y(_00558_));
 sky130_fd_sc_hd__nor2_2 _08492_ (.A(_00463_),
    .B(_00558_),
    .Y(_00559_));
 sky130_fd_sc_hd__nand2_2 _08493_ (.A(_00558_),
    .B(_00463_),
    .Y(_00560_));
 sky130_fd_sc_hd__and2b_1 _08494_ (.A_N(_00559_),
    .B(_00560_),
    .X(_00561_));
 sky130_fd_sc_hd__xnor2_2 _08495_ (.A(_00439_),
    .B(_00561_),
    .Y(_00562_));
 sky130_fd_sc_hd__o21ai_2 _08496_ (.A1(_04334_),
    .A2(_00348_),
    .B1(_04004_),
    .Y(_00564_));
 sky130_fd_sc_hd__and3_4 _08497_ (.A(_00412_),
    .B(_00562_),
    .C(_00564_),
    .X(_00565_));
 sky130_fd_sc_hd__a21oi_2 _08498_ (.A1(_00412_),
    .A2(_00564_),
    .B1(_00562_),
    .Y(_00566_));
 sky130_fd_sc_hd__nor2_2 _08499_ (.A(_00565_),
    .B(_00566_),
    .Y(_00567_));
 sky130_fd_sc_hd__inv_2 _08500_ (.A(_00371_),
    .Y(_00568_));
 sky130_fd_sc_hd__a22oi_4 _08501_ (.A1(_00350_),
    .A2(_00568_),
    .B1(_00372_),
    .B2(_00411_),
    .Y(_00569_));
 sky130_fd_sc_hd__xnor2_4 _08502_ (.A(_00567_),
    .B(_00569_),
    .Y(net77));
 sky130_fd_sc_hd__a21bo_1 _08503_ (.A1(_00417_),
    .A2(_00436_),
    .B1_N(_00437_),
    .X(_00570_));
 sky130_fd_sc_hd__buf_2 _08504_ (.A(net14),
    .X(_00571_));
 sky130_fd_sc_hd__clkbuf_4 _08505_ (.A(_00571_),
    .X(_00572_));
 sky130_fd_sc_hd__clkbuf_4 _08506_ (.A(_00572_),
    .X(_00574_));
 sky130_fd_sc_hd__clkbuf_4 _08507_ (.A(_00574_),
    .X(_00575_));
 sky130_fd_sc_hd__a22o_1 _08508_ (.A1(_02138_),
    .A2(_00415_),
    .B1(_00575_),
    .B2(_00333_),
    .X(_00576_));
 sky130_fd_sc_hd__and4_1 _08509_ (.A(_01744_),
    .B(_00311_),
    .C(_00413_),
    .D(_00571_),
    .X(_00577_));
 sky130_fd_sc_hd__inv_2 _08510_ (.A(_00577_),
    .Y(_00578_));
 sky130_fd_sc_hd__and2_1 _08511_ (.A(_00576_),
    .B(_00578_),
    .X(_00579_));
 sky130_fd_sc_hd__nand2_1 _08512_ (.A(_00421_),
    .B(_00427_),
    .Y(_00580_));
 sky130_fd_sc_hd__a22o_1 _08513_ (.A1(_01295_),
    .A2(_03894_),
    .B1(_03938_),
    .B2(_01405_),
    .X(_00581_));
 sky130_fd_sc_hd__nand4_1 _08514_ (.A(_01361_),
    .B(_01405_),
    .C(_03773_),
    .D(_03938_),
    .Y(_00582_));
 sky130_fd_sc_hd__o211a_1 _08515_ (.A1(_00422_),
    .A2(_00425_),
    .B1(_00581_),
    .C1(_00582_),
    .X(_00583_));
 sky130_fd_sc_hd__a211oi_1 _08516_ (.A1(_00581_),
    .A2(_00582_),
    .B1(_00422_),
    .C1(_00425_),
    .Y(_00585_));
 sky130_fd_sc_hd__nor2_1 _08517_ (.A(_00583_),
    .B(_00585_),
    .Y(_00586_));
 sky130_fd_sc_hd__xor2_2 _08518_ (.A(_00580_),
    .B(_00586_),
    .X(_00587_));
 sky130_fd_sc_hd__a21boi_2 _08519_ (.A1(_03982_),
    .A2(_00430_),
    .B1_N(_00429_),
    .Y(_00588_));
 sky130_fd_sc_hd__xor2_2 _08520_ (.A(_00587_),
    .B(net160),
    .X(_00589_));
 sky130_fd_sc_hd__a22o_1 _08521_ (.A1(_03059_),
    .A2(_00389_),
    .B1(_00393_),
    .B2(_02280_),
    .X(_00590_));
 sky130_fd_sc_hd__nand4_4 _08522_ (.A(_02007_),
    .B(_02040_),
    .C(_03707_),
    .D(_00392_),
    .Y(_00591_));
 sky130_fd_sc_hd__and2_1 _08523_ (.A(_00590_),
    .B(_00591_),
    .X(_00592_));
 sky130_fd_sc_hd__xor2_1 _08524_ (.A(_00589_),
    .B(_00592_),
    .X(_00593_));
 sky130_fd_sc_hd__xnor2_1 _08525_ (.A(_00579_),
    .B(_00593_),
    .Y(_00594_));
 sky130_fd_sc_hd__or2_4 _08526_ (.A(_00570_),
    .B(_00594_),
    .X(_00596_));
 sky130_fd_sc_hd__nand2_1 _08527_ (.A(_00570_),
    .B(_00594_),
    .Y(_00597_));
 sky130_fd_sc_hd__and2_2 _08528_ (.A(_00596_),
    .B(_00597_),
    .X(_00598_));
 sky130_fd_sc_hd__o21ai_1 _08529_ (.A1(_00454_),
    .A2(_00455_),
    .B1(_00461_),
    .Y(_00599_));
 sky130_fd_sc_hd__a32o_1 _08530_ (.A1(_00453_),
    .A2(_00460_),
    .A3(_00456_),
    .B1(_02467_),
    .B2(_00380_),
    .X(_00600_));
 sky130_fd_sc_hd__a22oi_1 _08531_ (.A1(_02259_),
    .A2(_00376_),
    .B1(_00379_),
    .B2(_02171_),
    .Y(_00601_));
 sky130_fd_sc_hd__and4_1 _08532_ (.A(_02105_),
    .B(_02149_),
    .C(_04037_),
    .D(_04048_),
    .X(_00602_));
 sky130_fd_sc_hd__or2_1 _08533_ (.A(_00601_),
    .B(_00602_),
    .X(_00603_));
 sky130_fd_sc_hd__clkbuf_4 _08534_ (.A(net46),
    .X(_00604_));
 sky130_fd_sc_hd__clkbuf_4 _08535_ (.A(_00604_),
    .X(_00605_));
 sky130_fd_sc_hd__clkbuf_4 _08536_ (.A(_00605_),
    .X(_00607_));
 sky130_fd_sc_hd__buf_4 _08537_ (.A(_00607_),
    .X(_00608_));
 sky130_fd_sc_hd__a22o_1 _08538_ (.A1(_02051_),
    .A2(_00458_),
    .B1(_00608_),
    .B2(_00442_),
    .X(_00609_));
 sky130_fd_sc_hd__nand4_1 _08539_ (.A(_00453_),
    .B(_02051_),
    .C(_00458_),
    .D(_00608_),
    .Y(_00610_));
 sky130_fd_sc_hd__a31oi_2 _08540_ (.A1(_04268_),
    .A2(_04026_),
    .A3(_00446_),
    .B1(_00445_),
    .Y(_00611_));
 sky130_fd_sc_hd__clkbuf_4 _08541_ (.A(_04103_),
    .X(_00612_));
 sky130_fd_sc_hd__clkbuf_4 _08542_ (.A(_04191_),
    .X(_00613_));
 sky130_fd_sc_hd__a22o_1 _08543_ (.A1(_01230_),
    .A2(_00612_),
    .B1(_00613_),
    .B2(_01284_),
    .X(_00614_));
 sky130_fd_sc_hd__nand4_1 _08544_ (.A(_01372_),
    .B(_04268_),
    .C(_00612_),
    .D(_00613_),
    .Y(_00615_));
 sky130_fd_sc_hd__nand2_1 _08545_ (.A(_00614_),
    .B(_00615_),
    .Y(_00616_));
 sky130_fd_sc_hd__xor2_1 _08546_ (.A(_00611_),
    .B(_00616_),
    .X(_00618_));
 sky130_fd_sc_hd__and3_1 _08547_ (.A(_00444_),
    .B(_00449_),
    .C(_00618_),
    .X(_00619_));
 sky130_fd_sc_hd__a21oi_1 _08548_ (.A1(_00444_),
    .A2(_00449_),
    .B1(_00618_),
    .Y(_00620_));
 sky130_fd_sc_hd__or2_1 _08549_ (.A(_00619_),
    .B(_00620_),
    .X(_00621_));
 sky130_fd_sc_hd__a21boi_2 _08550_ (.A1(_04312_),
    .A2(_00452_),
    .B1_N(_00451_),
    .Y(_00622_));
 sky130_fd_sc_hd__xor2_1 _08551_ (.A(_00621_),
    .B(_00622_),
    .X(_00623_));
 sky130_fd_sc_hd__a21oi_1 _08552_ (.A1(_00609_),
    .A2(_00610_),
    .B1(_00623_),
    .Y(_00624_));
 sky130_fd_sc_hd__and3_1 _08553_ (.A(_00623_),
    .B(_00609_),
    .C(_00610_),
    .X(_00625_));
 sky130_fd_sc_hd__nor2_1 _08554_ (.A(_00624_),
    .B(_00625_),
    .Y(_00626_));
 sky130_fd_sc_hd__xnor2_1 _08555_ (.A(_00603_),
    .B(_00626_),
    .Y(_00627_));
 sky130_fd_sc_hd__and3_1 _08556_ (.A(_00599_),
    .B(_00600_),
    .C(_00627_),
    .X(_00629_));
 sky130_fd_sc_hd__a21oi_1 _08557_ (.A1(_00599_),
    .A2(_00600_),
    .B1(_00627_),
    .Y(_00630_));
 sky130_fd_sc_hd__or2_1 _08558_ (.A(_00629_),
    .B(_00630_),
    .X(_00631_));
 sky130_fd_sc_hd__nand3_1 _08559_ (.A(_00410_),
    .B(_00544_),
    .C(_00542_),
    .Y(_00632_));
 sky130_fd_sc_hd__and2b_1 _08560_ (.A_N(_00542_),
    .B(_00545_),
    .X(_00633_));
 sky130_fd_sc_hd__a21o_1 _08561_ (.A1(_00527_),
    .A2(_00632_),
    .B1(_00633_),
    .X(_00634_));
 sky130_fd_sc_hd__buf_2 _08562_ (.A(_04917_),
    .X(_00635_));
 sky130_fd_sc_hd__clkbuf_4 _08563_ (.A(_00635_),
    .X(_00636_));
 sky130_fd_sc_hd__a22o_1 _08564_ (.A1(_00519_),
    .A2(_00636_),
    .B1(_00526_),
    .B2(_03554_),
    .X(_00637_));
 sky130_fd_sc_hd__and4_1 _08565_ (.A(_03554_),
    .B(_00508_),
    .C(_04917_),
    .D(_04939_),
    .X(_00638_));
 sky130_fd_sc_hd__inv_2 _08566_ (.A(_00638_),
    .Y(_00640_));
 sky130_fd_sc_hd__and2_1 _08567_ (.A(_00637_),
    .B(_00640_),
    .X(_00641_));
 sky130_fd_sc_hd__nand2_1 _08568_ (.A(_00531_),
    .B(_00536_),
    .Y(_00642_));
 sky130_fd_sc_hd__a31o_1 _08569_ (.A1(_03543_),
    .A2(_00294_),
    .A3(_00533_),
    .B1(_00532_),
    .X(_00643_));
 sky130_fd_sc_hd__a22oi_1 _08570_ (.A1(_06965_),
    .A2(_00293_),
    .B1(_00151_),
    .B2(_00263_),
    .Y(_00644_));
 sky130_fd_sc_hd__and4_1 _08571_ (.A(_06965_),
    .B(_06966_),
    .C(_00095_),
    .D(_00151_),
    .X(_00645_));
 sky130_fd_sc_hd__nor2_1 _08572_ (.A(_00644_),
    .B(_00645_),
    .Y(_00646_));
 sky130_fd_sc_hd__xnor2_1 _08573_ (.A(_00643_),
    .B(_00646_),
    .Y(_00647_));
 sky130_fd_sc_hd__nor2_1 _08574_ (.A(_00642_),
    .B(_00647_),
    .Y(_00648_));
 sky130_fd_sc_hd__and2_1 _08575_ (.A(_00642_),
    .B(_00647_),
    .X(_00649_));
 sky130_fd_sc_hd__nor2_1 _08576_ (.A(_00648_),
    .B(_00649_),
    .Y(_00651_));
 sky130_fd_sc_hd__o21ba_1 _08577_ (.A1(_00340_),
    .A2(_00539_),
    .B1_N(_00538_),
    .X(_00652_));
 sky130_fd_sc_hd__xnor2_1 _08578_ (.A(_00651_),
    .B(_00652_),
    .Y(_00653_));
 sky130_fd_sc_hd__buf_4 _08579_ (.A(_00004_),
    .X(_00654_));
 sky130_fd_sc_hd__a22o_1 _08580_ (.A1(_00399_),
    .A2(_00654_),
    .B1(_00543_),
    .B2(_03015_),
    .X(_00655_));
 sky130_fd_sc_hd__and3_1 _08581_ (.A(_00388_),
    .B(_02993_),
    .C(_06765_),
    .X(_00656_));
 sky130_fd_sc_hd__nand2_1 _08582_ (.A(_00543_),
    .B(_00656_),
    .Y(_00657_));
 sky130_fd_sc_hd__nand2_1 _08583_ (.A(_00655_),
    .B(_00657_),
    .Y(_00658_));
 sky130_fd_sc_hd__and2b_1 _08584_ (.A_N(_00653_),
    .B(_00658_),
    .X(_00659_));
 sky130_fd_sc_hd__and3_1 _08585_ (.A(_00653_),
    .B(_00655_),
    .C(_00657_),
    .X(_00660_));
 sky130_fd_sc_hd__nor2_1 _08586_ (.A(_00659_),
    .B(_00660_),
    .Y(_00662_));
 sky130_fd_sc_hd__xnor2_1 _08587_ (.A(_00641_),
    .B(_00662_),
    .Y(_00663_));
 sky130_fd_sc_hd__nor2_1 _08588_ (.A(_00634_),
    .B(_00663_),
    .Y(_00664_));
 sky130_fd_sc_hd__and2_1 _08589_ (.A(_00634_),
    .B(_00663_),
    .X(_00665_));
 sky130_fd_sc_hd__or2_2 _08590_ (.A(_00664_),
    .B(_00665_),
    .X(_00666_));
 sky130_fd_sc_hd__nor2_1 _08591_ (.A(_00493_),
    .B(_00523_),
    .Y(_00667_));
 sky130_fd_sc_hd__a21o_1 _08592_ (.A1(_00469_),
    .A2(_00492_),
    .B1(_00490_),
    .X(_00668_));
 sky130_fd_sc_hd__a31o_1 _08593_ (.A1(_06494_),
    .A2(_00004_),
    .A3(_00471_),
    .B1(_00472_),
    .X(_00669_));
 sky130_fd_sc_hd__buf_4 _08594_ (.A(_00258_),
    .X(_00670_));
 sky130_fd_sc_hd__a22oi_2 _08595_ (.A1(_06472_),
    .A2(_00257_),
    .B1(_00670_),
    .B2(_06483_),
    .Y(_00671_));
 sky130_fd_sc_hd__and4_1 _08596_ (.A(_06472_),
    .B(_06483_),
    .C(_00113_),
    .D(_00258_),
    .X(_00673_));
 sky130_fd_sc_hd__nor2_1 _08597_ (.A(_00671_),
    .B(_00673_),
    .Y(_00674_));
 sky130_fd_sc_hd__xor2_1 _08598_ (.A(_00669_),
    .B(_00674_),
    .X(_00675_));
 sky130_fd_sc_hd__and2_1 _08599_ (.A(_00479_),
    .B(_00675_),
    .X(_00676_));
 sky130_fd_sc_hd__nor2_1 _08600_ (.A(_00479_),
    .B(_00675_),
    .Y(_00677_));
 sky130_fd_sc_hd__or2_1 _08601_ (.A(_00676_),
    .B(_00677_),
    .X(_00678_));
 sky130_fd_sc_hd__and2b_1 _08602_ (.A_N(_00481_),
    .B(_00470_),
    .X(_00679_));
 sky130_fd_sc_hd__a21oi_1 _08603_ (.A1(_00280_),
    .A2(_00482_),
    .B1(_00679_),
    .Y(_00680_));
 sky130_fd_sc_hd__nor2_1 _08604_ (.A(_00678_),
    .B(_00680_),
    .Y(_00681_));
 sky130_fd_sc_hd__and2_1 _08605_ (.A(_00678_),
    .B(_00680_),
    .X(_00682_));
 sky130_fd_sc_hd__nor2_1 _08606_ (.A(_00681_),
    .B(_00682_),
    .Y(_00684_));
 sky130_fd_sc_hd__xnor2_2 _08607_ (.A(_00484_),
    .B(_00684_),
    .Y(_00685_));
 sky130_fd_sc_hd__xnor2_2 _08608_ (.A(_00668_),
    .B(_00685_),
    .Y(_00686_));
 sky130_fd_sc_hd__a21o_1 _08609_ (.A1(_00496_),
    .A2(_00522_),
    .B1(_00520_),
    .X(_00687_));
 sky130_fd_sc_hd__o21ba_1 _08610_ (.A1(_00316_),
    .A2(_00510_),
    .B1_N(_00509_),
    .X(_00688_));
 sky130_fd_sc_hd__a22oi_1 _08611_ (.A1(_06428_),
    .A2(_00144_),
    .B1(_00310_),
    .B2(_06450_),
    .Y(_00689_));
 sky130_fd_sc_hd__and4_1 _08612_ (.A(_06428_),
    .B(_06439_),
    .C(_00144_),
    .D(_00298_),
    .X(_00690_));
 sky130_fd_sc_hd__nor2_1 _08613_ (.A(_00689_),
    .B(_00690_),
    .Y(_00691_));
 sky130_fd_sc_hd__o21a_1 _08614_ (.A1(_00500_),
    .A2(_00502_),
    .B1(_00691_),
    .X(_00692_));
 sky130_fd_sc_hd__nor3_1 _08615_ (.A(_00500_),
    .B(_00502_),
    .C(_00691_),
    .Y(_00693_));
 sky130_fd_sc_hd__nor2_1 _08616_ (.A(_00692_),
    .B(_00693_),
    .Y(_00695_));
 sky130_fd_sc_hd__and2_1 _08617_ (.A(_00505_),
    .B(_00695_),
    .X(_00696_));
 sky130_fd_sc_hd__nor2_1 _08618_ (.A(_00505_),
    .B(_00695_),
    .Y(_00697_));
 sky130_fd_sc_hd__nor2_1 _08619_ (.A(_00696_),
    .B(_00697_),
    .Y(_00698_));
 sky130_fd_sc_hd__and2b_1 _08620_ (.A_N(_00688_),
    .B(_00698_),
    .X(_00699_));
 sky130_fd_sc_hd__and2b_1 _08621_ (.A_N(_00698_),
    .B(_00688_),
    .X(_00700_));
 sky130_fd_sc_hd__nor2_2 _08622_ (.A(_00699_),
    .B(_00700_),
    .Y(_00701_));
 sky130_fd_sc_hd__xnor2_4 _08623_ (.A(_00513_),
    .B(_00701_),
    .Y(_00702_));
 sky130_fd_sc_hd__xnor2_4 _08624_ (.A(_00687_),
    .B(_00702_),
    .Y(_00703_));
 sky130_fd_sc_hd__xor2_2 _08625_ (.A(_00686_),
    .B(_00703_),
    .X(_00704_));
 sky130_fd_sc_hd__xor2_1 _08626_ (.A(_00667_),
    .B(_00704_),
    .X(_00706_));
 sky130_fd_sc_hd__xnor2_2 _08627_ (.A(_00666_),
    .B(_00706_),
    .Y(_00707_));
 sky130_fd_sc_hd__a21o_1 _08628_ (.A1(_00466_),
    .A2(_00524_),
    .B1(_00547_),
    .X(_00708_));
 sky130_fd_sc_hd__o21a_1 _08629_ (.A1(_00466_),
    .A2(_00524_),
    .B1(_00708_),
    .X(_00709_));
 sky130_fd_sc_hd__xnor2_2 _08630_ (.A(_00707_),
    .B(_00709_),
    .Y(_00710_));
 sky130_fd_sc_hd__inv_2 _08631_ (.A(_00550_),
    .Y(_00711_));
 sky130_fd_sc_hd__and3b_1 _08632_ (.A_N(_00551_),
    .B(_00347_),
    .C(_00711_),
    .X(_00712_));
 sky130_fd_sc_hd__a21oi_1 _08633_ (.A1(_00555_),
    .A2(_00711_),
    .B1(_00551_),
    .Y(_00713_));
 sky130_fd_sc_hd__a21oi_1 _08634_ (.A1(_00251_),
    .A2(_00712_),
    .B1(_00713_),
    .Y(_00714_));
 sky130_fd_sc_hd__xnor2_2 _08635_ (.A(_00710_),
    .B(_00714_),
    .Y(_00715_));
 sky130_fd_sc_hd__xnor2_1 _08636_ (.A(_00631_),
    .B(_00715_),
    .Y(_00717_));
 sky130_fd_sc_hd__xnor2_2 _08637_ (.A(_00598_),
    .B(_00717_),
    .Y(_00718_));
 sky130_fd_sc_hd__a21oi_2 _08638_ (.A1(_00439_),
    .A2(_00560_),
    .B1(_00559_),
    .Y(_00719_));
 sky130_fd_sc_hd__xnor2_1 _08639_ (.A(_00718_),
    .B(_00719_),
    .Y(_00720_));
 sky130_fd_sc_hd__or4_4 _08640_ (.A(_00565_),
    .B(_00566_),
    .C(_00569_),
    .D(_00720_),
    .X(_00721_));
 sky130_fd_sc_hd__xor2_1 _08641_ (.A(_00718_),
    .B(_00719_),
    .X(_00722_));
 sky130_fd_sc_hd__xnor2_1 _08642_ (.A(_00565_),
    .B(_00722_),
    .Y(_00723_));
 sky130_fd_sc_hd__o31ai_1 _08643_ (.A1(_00565_),
    .A2(_00566_),
    .A3(_00569_),
    .B1(_00723_),
    .Y(_00724_));
 sky130_fd_sc_hd__and2_4 _08644_ (.A(_00721_),
    .B(_00724_),
    .X(_00725_));
 sky130_fd_sc_hd__clkbuf_1 _08645_ (.A(_00725_),
    .X(net78));
 sky130_fd_sc_hd__and2_2 _08646_ (.A(_00718_),
    .B(_00719_),
    .X(_00727_));
 sky130_fd_sc_hd__o21a_1 _08647_ (.A1(_00589_),
    .A2(_00592_),
    .B1(_00579_),
    .X(_00728_));
 sky130_fd_sc_hd__a31o_2 _08648_ (.A1(_00589_),
    .A2(_00590_),
    .A3(_00591_),
    .B1(_00728_),
    .X(_00729_));
 sky130_fd_sc_hd__buf_2 _08649_ (.A(net14),
    .X(_00730_));
 sky130_fd_sc_hd__and4_1 _08650_ (.A(_04510_),
    .B(_00661_),
    .C(net13),
    .D(_00730_),
    .X(_00731_));
 sky130_fd_sc_hd__a22o_1 _08651_ (.A1(_01394_),
    .A2(net13),
    .B1(_00730_),
    .B2(_01470_),
    .X(_00732_));
 sky130_fd_sc_hd__or2b_1 _08652_ (.A(_00731_),
    .B_N(_00732_),
    .X(_00733_));
 sky130_fd_sc_hd__clkbuf_4 _08653_ (.A(net15),
    .X(_00734_));
 sky130_fd_sc_hd__nand2_1 _08654_ (.A(_00311_),
    .B(_00734_),
    .Y(_00735_));
 sky130_fd_sc_hd__xnor2_1 _08655_ (.A(_00733_),
    .B(_00735_),
    .Y(_00736_));
 sky130_fd_sc_hd__or2_1 _08656_ (.A(_00578_),
    .B(_00736_),
    .X(_00738_));
 sky130_fd_sc_hd__nand2_1 _08657_ (.A(_00578_),
    .B(_00736_),
    .Y(_00739_));
 sky130_fd_sc_hd__and2_2 _08658_ (.A(_00738_),
    .B(_00739_),
    .X(_00740_));
 sky130_fd_sc_hd__clkbuf_4 _08659_ (.A(_03938_),
    .X(_00741_));
 sky130_fd_sc_hd__buf_4 _08660_ (.A(_03773_),
    .X(_00742_));
 sky130_fd_sc_hd__nand2_1 _08661_ (.A(_00159_),
    .B(_00742_),
    .Y(_00743_));
 sky130_fd_sc_hd__and4_1 _08662_ (.A(_00157_),
    .B(_00741_),
    .C(_00743_),
    .D(_00583_),
    .X(_00744_));
 sky130_fd_sc_hd__buf_4 _08663_ (.A(_00741_),
    .X(_00745_));
 sky130_fd_sc_hd__a31o_1 _08664_ (.A1(_00157_),
    .A2(_00745_),
    .A3(_00743_),
    .B1(_00583_),
    .X(_00746_));
 sky130_fd_sc_hd__and2b_1 _08665_ (.A_N(_00744_),
    .B(_00746_),
    .X(_00747_));
 sky130_fd_sc_hd__and3_1 _08666_ (.A(_00421_),
    .B(_00427_),
    .C(_00586_),
    .X(_00749_));
 sky130_fd_sc_hd__o21bai_2 _08667_ (.A1(_00587_),
    .A2(_00588_),
    .B1_N(_00749_),
    .Y(_00750_));
 sky130_fd_sc_hd__xnor2_2 _08668_ (.A(_00747_),
    .B(_00750_),
    .Y(_00751_));
 sky130_fd_sc_hd__and4_1 _08669_ (.A(_05731_),
    .B(net60),
    .C(net8),
    .D(net9),
    .X(_00752_));
 sky130_fd_sc_hd__a22o_1 _08670_ (.A1(_05731_),
    .A2(net8),
    .B1(_03718_),
    .B2(_01000_),
    .X(_00753_));
 sky130_fd_sc_hd__or2b_1 _08671_ (.A(_00752_),
    .B_N(_00753_),
    .X(_00754_));
 sky130_fd_sc_hd__buf_4 _08672_ (.A(_03894_),
    .X(_00755_));
 sky130_fd_sc_hd__nand2_1 _08673_ (.A(_02029_),
    .B(_00755_),
    .Y(_00756_));
 sky130_fd_sc_hd__xnor2_1 _08674_ (.A(_00754_),
    .B(_00756_),
    .Y(_00757_));
 sky130_fd_sc_hd__nor2_1 _08675_ (.A(_00591_),
    .B(_00757_),
    .Y(_00758_));
 sky130_fd_sc_hd__and2_1 _08676_ (.A(_00591_),
    .B(_00757_),
    .X(_00760_));
 sky130_fd_sc_hd__or2_2 _08677_ (.A(_00758_),
    .B(_00760_),
    .X(_00761_));
 sky130_fd_sc_hd__xnor2_2 _08678_ (.A(_00751_),
    .B(_00761_),
    .Y(_00762_));
 sky130_fd_sc_hd__xnor2_4 _08679_ (.A(_00740_),
    .B(_00762_),
    .Y(_00763_));
 sky130_fd_sc_hd__xnor2_4 _08680_ (.A(_00729_),
    .B(_00763_),
    .Y(_00764_));
 sky130_fd_sc_hd__xnor2_4 _08681_ (.A(_00596_),
    .B(_00764_),
    .Y(_00765_));
 sky130_fd_sc_hd__o21ba_1 _08682_ (.A1(_00603_),
    .A2(_00624_),
    .B1_N(_00625_),
    .X(_00766_));
 sky130_fd_sc_hd__and4_1 _08683_ (.A(_00563_),
    .B(_00639_),
    .C(_04015_),
    .D(_04103_),
    .X(_00767_));
 sky130_fd_sc_hd__a22o_1 _08684_ (.A1(_00639_),
    .A2(_04015_),
    .B1(_04103_),
    .B2(_00563_),
    .X(_00768_));
 sky130_fd_sc_hd__and2b_1 _08685_ (.A_N(_00767_),
    .B(_00768_),
    .X(_00769_));
 sky130_fd_sc_hd__nand2_1 _08686_ (.A(_05577_),
    .B(_04048_),
    .Y(_00771_));
 sky130_fd_sc_hd__xnor2_1 _08687_ (.A(_00769_),
    .B(_00771_),
    .Y(_00772_));
 sky130_fd_sc_hd__and2_1 _08688_ (.A(_00602_),
    .B(_00772_),
    .X(_00773_));
 sky130_fd_sc_hd__nor2_1 _08689_ (.A(_00602_),
    .B(_00772_),
    .Y(_00774_));
 sky130_fd_sc_hd__nor2_1 _08690_ (.A(_00773_),
    .B(_00774_),
    .Y(_00775_));
 sky130_fd_sc_hd__nor2_1 _08691_ (.A(_00611_),
    .B(_00616_),
    .Y(_00776_));
 sky130_fd_sc_hd__buf_2 _08692_ (.A(net43),
    .X(_00777_));
 sky130_fd_sc_hd__clkbuf_4 _08693_ (.A(_00777_),
    .X(_00778_));
 sky130_fd_sc_hd__clkbuf_4 _08694_ (.A(_00778_),
    .X(_00779_));
 sky130_fd_sc_hd__buf_2 _08695_ (.A(_04180_),
    .X(_00780_));
 sky130_fd_sc_hd__clkbuf_4 _08696_ (.A(_00780_),
    .X(_00782_));
 sky130_fd_sc_hd__buf_2 _08697_ (.A(_00782_),
    .X(_00783_));
 sky130_fd_sc_hd__clkbuf_4 _08698_ (.A(_00783_),
    .X(_00784_));
 sky130_fd_sc_hd__nand2_1 _08699_ (.A(_01383_),
    .B(_00784_),
    .Y(_00785_));
 sky130_fd_sc_hd__and3_2 _08700_ (.A(_01350_),
    .B(_00779_),
    .C(_00785_),
    .X(_00786_));
 sky130_fd_sc_hd__xor2_2 _08701_ (.A(_00776_),
    .B(_00786_),
    .X(_00787_));
 sky130_fd_sc_hd__o21bai_2 _08702_ (.A1(_00621_),
    .A2(_00622_),
    .B1_N(_00619_),
    .Y(_00788_));
 sky130_fd_sc_hd__xnor2_2 _08703_ (.A(_00787_),
    .B(_00788_),
    .Y(_00789_));
 sky130_fd_sc_hd__and4_1 _08704_ (.A(_00442_),
    .B(_00989_),
    .C(net45),
    .D(_00604_),
    .X(_00790_));
 sky130_fd_sc_hd__and4_1 _08705_ (.A(_00431_),
    .B(_04169_),
    .C(net46),
    .D(net47),
    .X(_00791_));
 sky130_fd_sc_hd__a22o_1 _08706_ (.A1(_03587_),
    .A2(net46),
    .B1(net47),
    .B2(_00431_),
    .X(_00793_));
 sky130_fd_sc_hd__and2b_1 _08707_ (.A_N(_00791_),
    .B(_00793_),
    .X(_00794_));
 sky130_fd_sc_hd__nand2_1 _08708_ (.A(_04081_),
    .B(net45),
    .Y(_00795_));
 sky130_fd_sc_hd__xnor2_1 _08709_ (.A(_00794_),
    .B(_00795_),
    .Y(_00796_));
 sky130_fd_sc_hd__and2_1 _08710_ (.A(_00790_),
    .B(_00796_),
    .X(_00797_));
 sky130_fd_sc_hd__nor2_1 _08711_ (.A(_00790_),
    .B(_00796_),
    .Y(_00798_));
 sky130_fd_sc_hd__or2_1 _08712_ (.A(_00797_),
    .B(_00798_),
    .X(_00799_));
 sky130_fd_sc_hd__xnor2_1 _08713_ (.A(_00789_),
    .B(_00799_),
    .Y(_00800_));
 sky130_fd_sc_hd__xnor2_1 _08714_ (.A(_00775_),
    .B(_00800_),
    .Y(_00801_));
 sky130_fd_sc_hd__xnor2_1 _08715_ (.A(_00766_),
    .B(_00801_),
    .Y(_00802_));
 sky130_fd_sc_hd__xnor2_1 _08716_ (.A(_00629_),
    .B(_00802_),
    .Y(_00804_));
 sky130_fd_sc_hd__or2b_1 _08717_ (.A(_00653_),
    .B_N(_00658_),
    .X(_00805_));
 sky130_fd_sc_hd__a21oi_1 _08718_ (.A1(_00641_),
    .A2(_00805_),
    .B1(_00660_),
    .Y(_00806_));
 sky130_fd_sc_hd__and4_1 _08719_ (.A(_03532_),
    .B(_00121_),
    .C(_04895_),
    .D(_04873_),
    .X(_00807_));
 sky130_fd_sc_hd__a22o_1 _08720_ (.A1(_03532_),
    .A2(_04895_),
    .B1(_04873_),
    .B2(_00121_),
    .X(_00808_));
 sky130_fd_sc_hd__and4b_1 _08721_ (.A_N(_00807_),
    .B(_00808_),
    .C(_00497_),
    .D(_00142_),
    .X(_00809_));
 sky130_fd_sc_hd__inv_2 _08722_ (.A(_00808_),
    .Y(_00810_));
 sky130_fd_sc_hd__o2bb2a_1 _08723_ (.A1_N(_00508_),
    .A2_N(_00144_),
    .B1(_00807_),
    .B2(_00810_),
    .X(_00811_));
 sky130_fd_sc_hd__or2_1 _08724_ (.A(_00809_),
    .B(_00811_),
    .X(_00812_));
 sky130_fd_sc_hd__or2_1 _08725_ (.A(_00640_),
    .B(_00812_),
    .X(_00813_));
 sky130_fd_sc_hd__nand2_1 _08726_ (.A(_00640_),
    .B(_00812_),
    .Y(_00815_));
 sky130_fd_sc_hd__nand2_1 _08727_ (.A(_00813_),
    .B(_00815_),
    .Y(_00816_));
 sky130_fd_sc_hd__and2_1 _08728_ (.A(_00643_),
    .B(_00646_),
    .X(_00817_));
 sky130_fd_sc_hd__clkbuf_4 _08729_ (.A(_00294_),
    .X(_00818_));
 sky130_fd_sc_hd__clkbuf_4 _08730_ (.A(_00293_),
    .X(_00819_));
 sky130_fd_sc_hd__nand2_1 _08731_ (.A(_00263_),
    .B(_00819_),
    .Y(_00820_));
 sky130_fd_sc_hd__and3_1 _08732_ (.A(_00262_),
    .B(_00818_),
    .C(_00820_),
    .X(_00821_));
 sky130_fd_sc_hd__xor2_1 _08733_ (.A(_00817_),
    .B(_00821_),
    .X(_00822_));
 sky130_fd_sc_hd__o21bai_1 _08734_ (.A1(_00649_),
    .A2(_00652_),
    .B1_N(_00648_),
    .Y(_00823_));
 sky130_fd_sc_hd__xnor2_1 _08735_ (.A(_00822_),
    .B(_00823_),
    .Y(_00824_));
 sky130_fd_sc_hd__a22o_1 _08736_ (.A1(_00377_),
    .A2(_00114_),
    .B1(_06765_),
    .B2(_02993_),
    .X(_00826_));
 sky130_fd_sc_hd__a21bo_1 _08737_ (.A1(_00258_),
    .A2(_00656_),
    .B1_N(_00826_),
    .X(_00827_));
 sky130_fd_sc_hd__nand2_1 _08738_ (.A(_06885_),
    .B(_00293_),
    .Y(_00828_));
 sky130_fd_sc_hd__xor2_1 _08739_ (.A(_00827_),
    .B(_00828_),
    .X(_00829_));
 sky130_fd_sc_hd__and3_1 _08740_ (.A(_07004_),
    .B(_00656_),
    .C(_00829_),
    .X(_00830_));
 sky130_fd_sc_hd__a21oi_1 _08741_ (.A1(_00543_),
    .A2(_00656_),
    .B1(_00829_),
    .Y(_00831_));
 sky130_fd_sc_hd__or2_1 _08742_ (.A(_00830_),
    .B(_00831_),
    .X(_00832_));
 sky130_fd_sc_hd__nand2_1 _08743_ (.A(_00824_),
    .B(_00832_),
    .Y(_00833_));
 sky130_fd_sc_hd__or2_1 _08744_ (.A(_00824_),
    .B(_00832_),
    .X(_00834_));
 sky130_fd_sc_hd__nand2_1 _08745_ (.A(_00833_),
    .B(_00834_),
    .Y(_00835_));
 sky130_fd_sc_hd__xor2_1 _08746_ (.A(_00816_),
    .B(_00835_),
    .X(_00837_));
 sky130_fd_sc_hd__xnor2_1 _08747_ (.A(_00806_),
    .B(_00837_),
    .Y(_00838_));
 sky130_fd_sc_hd__nand2_1 _08748_ (.A(_00664_),
    .B(_00838_),
    .Y(_00839_));
 sky130_fd_sc_hd__or2_1 _08749_ (.A(_00664_),
    .B(_00838_),
    .X(_00840_));
 sky130_fd_sc_hd__and2_1 _08750_ (.A(_00839_),
    .B(_00840_),
    .X(_00841_));
 sky130_fd_sc_hd__nand2_1 _08751_ (.A(_00686_),
    .B(_00703_),
    .Y(_00842_));
 sky130_fd_sc_hd__clkbuf_4 _08752_ (.A(_00257_),
    .X(_00843_));
 sky130_fd_sc_hd__buf_4 _08753_ (.A(_00670_),
    .X(_00844_));
 sky130_fd_sc_hd__nand2_1 _08754_ (.A(_06937_),
    .B(_00844_),
    .Y(_00845_));
 sky130_fd_sc_hd__and3_1 _08755_ (.A(_06637_),
    .B(_00843_),
    .C(_00845_),
    .X(_00846_));
 sky130_fd_sc_hd__and3_1 _08756_ (.A(_00669_),
    .B(_00674_),
    .C(_00846_),
    .X(_00848_));
 sky130_fd_sc_hd__a21oi_1 _08757_ (.A1(_00669_),
    .A2(_00674_),
    .B1(_00846_),
    .Y(_00849_));
 sky130_fd_sc_hd__nor2_1 _08758_ (.A(_00848_),
    .B(_00849_),
    .Y(_00850_));
 sky130_fd_sc_hd__nor3_1 _08759_ (.A(_00676_),
    .B(_00681_),
    .C(_00850_),
    .Y(_00851_));
 sky130_fd_sc_hd__o21a_1 _08760_ (.A1(_00676_),
    .A2(_00681_),
    .B1(_00850_),
    .X(_00852_));
 sky130_fd_sc_hd__nor2_2 _08761_ (.A(_00851_),
    .B(_00852_),
    .Y(_00853_));
 sky130_fd_sc_hd__inv_2 _08762_ (.A(_00685_),
    .Y(_00854_));
 sky130_fd_sc_hd__o21a_1 _08763_ (.A1(_00484_),
    .A2(_00490_),
    .B1(_00684_),
    .X(_00855_));
 sky130_fd_sc_hd__a31o_1 _08764_ (.A1(_00469_),
    .A2(_00492_),
    .A3(_00854_),
    .B1(_00855_),
    .X(_00856_));
 sky130_fd_sc_hd__xor2_2 _08765_ (.A(_00853_),
    .B(_00856_),
    .X(_00857_));
 sky130_fd_sc_hd__clkbuf_4 _08766_ (.A(_00310_),
    .X(_00859_));
 sky130_fd_sc_hd__and3_1 _08767_ (.A(_06626_),
    .B(_00859_),
    .C(_00498_),
    .X(_00860_));
 sky130_fd_sc_hd__and2_1 _08768_ (.A(_00692_),
    .B(_00860_),
    .X(_00861_));
 sky130_fd_sc_hd__nor2_1 _08769_ (.A(_00692_),
    .B(_00860_),
    .Y(_00862_));
 sky130_fd_sc_hd__nor2_1 _08770_ (.A(_00861_),
    .B(_00862_),
    .Y(_00863_));
 sky130_fd_sc_hd__nor3_1 _08771_ (.A(_00696_),
    .B(_00699_),
    .C(_00863_),
    .Y(_00864_));
 sky130_fd_sc_hd__o21a_1 _08772_ (.A1(_00696_),
    .A2(_00699_),
    .B1(_00863_),
    .X(_00865_));
 sky130_fd_sc_hd__nor2_2 _08773_ (.A(_00864_),
    .B(_00865_),
    .Y(_00866_));
 sky130_fd_sc_hd__inv_2 _08774_ (.A(_00702_),
    .Y(_00867_));
 sky130_fd_sc_hd__o21a_1 _08775_ (.A1(_00513_),
    .A2(_00520_),
    .B1(_00701_),
    .X(_00868_));
 sky130_fd_sc_hd__a31oi_4 _08776_ (.A1(_00496_),
    .A2(_00522_),
    .A3(_00867_),
    .B1(_00868_),
    .Y(_00870_));
 sky130_fd_sc_hd__xnor2_4 _08777_ (.A(_00866_),
    .B(_00870_),
    .Y(_00871_));
 sky130_fd_sc_hd__xnor2_2 _08778_ (.A(_00857_),
    .B(_00871_),
    .Y(_00872_));
 sky130_fd_sc_hd__xnor2_1 _08779_ (.A(_00842_),
    .B(_00872_),
    .Y(_00873_));
 sky130_fd_sc_hd__xnor2_2 _08780_ (.A(_00841_),
    .B(_00873_),
    .Y(_00874_));
 sky130_fd_sc_hd__a21boi_1 _08781_ (.A1(_00667_),
    .A2(_00704_),
    .B1_N(_00666_),
    .Y(_00875_));
 sky130_fd_sc_hd__o21ba_1 _08782_ (.A1(_00667_),
    .A2(_00704_),
    .B1_N(_00875_),
    .X(_00876_));
 sky130_fd_sc_hd__xnor2_2 _08783_ (.A(_00874_),
    .B(_00876_),
    .Y(_00877_));
 sky130_fd_sc_hd__or2_1 _08784_ (.A(_00553_),
    .B(_00710_),
    .X(_00878_));
 sky130_fd_sc_hd__or3_1 _08785_ (.A(_00553_),
    .B(_00556_),
    .C(_00710_),
    .X(_00879_));
 sky130_fd_sc_hd__nand2_1 _08786_ (.A(_00707_),
    .B(_00709_),
    .Y(_00881_));
 sky130_fd_sc_hd__nor2_1 _08787_ (.A(_00707_),
    .B(_00709_),
    .Y(_00882_));
 sky130_fd_sc_hd__a21o_1 _08788_ (.A1(_00711_),
    .A2(_00881_),
    .B1(_00882_),
    .X(_00883_));
 sky130_fd_sc_hd__o311a_4 _08789_ (.A1(_00367_),
    .A2(_00554_),
    .A3(_00878_),
    .B1(_00879_),
    .C1(_00883_),
    .X(_00884_));
 sky130_fd_sc_hd__xnor2_1 _08790_ (.A(_00877_),
    .B(_00884_),
    .Y(_00885_));
 sky130_fd_sc_hd__and2_1 _08791_ (.A(_00804_),
    .B(_00885_),
    .X(_00886_));
 sky130_fd_sc_hd__or2_1 _08792_ (.A(_00804_),
    .B(_00885_),
    .X(_00887_));
 sky130_fd_sc_hd__and2b_1 _08793_ (.A_N(_00886_),
    .B(_00887_),
    .X(_00888_));
 sky130_fd_sc_hd__xnor2_2 _08794_ (.A(_00765_),
    .B(_00888_),
    .Y(_00889_));
 sky130_fd_sc_hd__o21bai_1 _08795_ (.A1(_00631_),
    .A2(_00715_),
    .B1_N(_00598_),
    .Y(_00890_));
 sky130_fd_sc_hd__a21bo_1 _08796_ (.A1(_00631_),
    .A2(_00715_),
    .B1_N(_00890_),
    .X(_00892_));
 sky130_fd_sc_hd__xnor2_2 _08797_ (.A(_00889_),
    .B(_00892_),
    .Y(_00893_));
 sky130_fd_sc_hd__xnor2_2 _08798_ (.A(_00727_),
    .B(_00893_),
    .Y(_00894_));
 sky130_fd_sc_hd__nand3_1 _08799_ (.A(_00412_),
    .B(_00562_),
    .C(_00564_),
    .Y(_00895_));
 sky130_fd_sc_hd__a211o_2 _08800_ (.A1(_00895_),
    .A2(_00569_),
    .B1(_00720_),
    .C1(_00566_),
    .X(_00896_));
 sky130_fd_sc_hd__xor2_2 _08801_ (.A(_00894_),
    .B(_00896_),
    .X(net79));
 sky130_fd_sc_hd__a21o_1 _08802_ (.A1(_00565_),
    .A2(_00722_),
    .B1(_00727_),
    .X(_00897_));
 sky130_fd_sc_hd__o2bb2a_4 _08803_ (.A1_N(_00893_),
    .A2_N(_00897_),
    .B1(_00894_),
    .B2(_00721_),
    .X(_00898_));
 sky130_fd_sc_hd__or2b_4 _08804_ (.A(_00889_),
    .B_N(_00892_),
    .X(_00899_));
 sky130_fd_sc_hd__and4_1 _08805_ (.A(_03850_),
    .B(_04510_),
    .C(net13),
    .D(_00730_),
    .X(_00900_));
 sky130_fd_sc_hd__a22o_1 _08806_ (.A1(_03850_),
    .A2(net13),
    .B1(_00730_),
    .B2(_01394_),
    .X(_00902_));
 sky130_fd_sc_hd__and2b_1 _08807_ (.A_N(_00900_),
    .B(_00902_),
    .X(_00903_));
 sky130_fd_sc_hd__nand2_1 _08808_ (.A(_02127_),
    .B(_00734_),
    .Y(_00904_));
 sky130_fd_sc_hd__xnor2_1 _08809_ (.A(_00903_),
    .B(_00904_),
    .Y(_00905_));
 sky130_fd_sc_hd__a31o_1 _08810_ (.A1(_00300_),
    .A2(net15),
    .A3(_00732_),
    .B1(_00731_),
    .X(_00906_));
 sky130_fd_sc_hd__and2_1 _08811_ (.A(_00300_),
    .B(net16),
    .X(_00907_));
 sky130_fd_sc_hd__xor2_1 _08812_ (.A(_00906_),
    .B(_00907_),
    .X(_00908_));
 sky130_fd_sc_hd__xnor2_1 _08813_ (.A(_00905_),
    .B(_00908_),
    .Y(_00909_));
 sky130_fd_sc_hd__nor2_1 _08814_ (.A(_00738_),
    .B(_00909_),
    .Y(_00910_));
 sky130_fd_sc_hd__and2_1 _08815_ (.A(_00738_),
    .B(_00909_),
    .X(_00911_));
 sky130_fd_sc_hd__or2_2 _08816_ (.A(_00910_),
    .B(_00911_),
    .X(_00913_));
 sky130_fd_sc_hd__clkbuf_4 _08817_ (.A(_00742_),
    .X(_00914_));
 sky130_fd_sc_hd__clkbuf_4 _08818_ (.A(_00914_),
    .X(_00915_));
 sky130_fd_sc_hd__clkbuf_4 _08819_ (.A(_00741_),
    .X(_00916_));
 sky130_fd_sc_hd__and4_1 _08820_ (.A(_00157_),
    .B(_00159_),
    .C(_00915_),
    .D(_00916_),
    .X(_00917_));
 sky130_fd_sc_hd__and2_1 _08821_ (.A(_00747_),
    .B(_00750_),
    .X(_00918_));
 sky130_fd_sc_hd__and4_1 _08822_ (.A(_01044_),
    .B(_05731_),
    .C(net8),
    .D(net9),
    .X(_00919_));
 sky130_fd_sc_hd__a22o_1 _08823_ (.A1(_01044_),
    .A2(net8),
    .B1(_03718_),
    .B2(_05731_),
    .X(_00920_));
 sky130_fd_sc_hd__and2b_1 _08824_ (.A_N(_00919_),
    .B(_00920_),
    .X(_00921_));
 sky130_fd_sc_hd__nand2_1 _08825_ (.A(_01996_),
    .B(_03762_),
    .Y(_00922_));
 sky130_fd_sc_hd__xnor2_1 _08826_ (.A(_00921_),
    .B(_00922_),
    .Y(_00924_));
 sky130_fd_sc_hd__a31o_1 _08827_ (.A1(_00901_),
    .A2(_03762_),
    .A3(_00753_),
    .B1(_00752_),
    .X(_00925_));
 sky130_fd_sc_hd__and2_1 _08828_ (.A(_00901_),
    .B(net11),
    .X(_00926_));
 sky130_fd_sc_hd__xor2_1 _08829_ (.A(_00925_),
    .B(_00926_),
    .X(_00927_));
 sky130_fd_sc_hd__xnor2_1 _08830_ (.A(_00924_),
    .B(_00927_),
    .Y(_00928_));
 sky130_fd_sc_hd__nor3_1 _08831_ (.A(_00591_),
    .B(_00757_),
    .C(_00928_),
    .Y(_00929_));
 sky130_fd_sc_hd__and2b_1 _08832_ (.A_N(_00758_),
    .B(_00928_),
    .X(_00930_));
 sky130_fd_sc_hd__nor2_1 _08833_ (.A(_00929_),
    .B(_00930_),
    .Y(_00931_));
 sky130_fd_sc_hd__or4_1 _08834_ (.A(_00917_),
    .B(_00744_),
    .C(_00918_),
    .D(_00931_),
    .X(_00932_));
 sky130_fd_sc_hd__o31ai_2 _08835_ (.A1(_00917_),
    .A2(_00744_),
    .A3(_00918_),
    .B1(_00931_),
    .Y(_00933_));
 sky130_fd_sc_hd__nand2_2 _08836_ (.A(_00932_),
    .B(_00933_),
    .Y(_00935_));
 sky130_fd_sc_hd__xor2_4 _08837_ (.A(_00913_),
    .B(_00935_),
    .X(_00936_));
 sky130_fd_sc_hd__nor2_1 _08838_ (.A(_00751_),
    .B(_00761_),
    .Y(_00937_));
 sky130_fd_sc_hd__nand2_1 _08839_ (.A(_00751_),
    .B(_00761_),
    .Y(_00938_));
 sky130_fd_sc_hd__o21ai_2 _08840_ (.A1(_00740_),
    .A2(_00937_),
    .B1(_00938_),
    .Y(_00939_));
 sky130_fd_sc_hd__xnor2_4 _08841_ (.A(_00936_),
    .B(_00939_),
    .Y(_00940_));
 sky130_fd_sc_hd__nand2_1 _08842_ (.A(_00729_),
    .B(_00763_),
    .Y(_00941_));
 sky130_fd_sc_hd__o21ai_4 _08843_ (.A1(_00596_),
    .A2(_00764_),
    .B1(_00941_),
    .Y(_00942_));
 sky130_fd_sc_hd__xnor2_4 _08844_ (.A(_00940_),
    .B(_00942_),
    .Y(_00943_));
 sky130_fd_sc_hd__and4_1 _08845_ (.A(_00563_),
    .B(_00639_),
    .C(_04180_),
    .D(_04191_),
    .X(_00944_));
 sky130_fd_sc_hd__a22o_1 _08846_ (.A1(_05742_),
    .A2(_04103_),
    .B1(_04191_),
    .B2(_00563_),
    .X(_00946_));
 sky130_fd_sc_hd__or2b_1 _08847_ (.A(_00944_),
    .B_N(_00946_),
    .X(_00947_));
 sky130_fd_sc_hd__nand2_1 _08848_ (.A(_05577_),
    .B(_04026_),
    .Y(_00948_));
 sky130_fd_sc_hd__xnor2_1 _08849_ (.A(_00947_),
    .B(_00948_),
    .Y(_00949_));
 sky130_fd_sc_hd__a31o_1 _08850_ (.A1(_02664_),
    .A2(net40),
    .A3(_00768_),
    .B1(_00767_),
    .X(_00950_));
 sky130_fd_sc_hd__and2_1 _08851_ (.A(_03268_),
    .B(net40),
    .X(_00951_));
 sky130_fd_sc_hd__xnor2_1 _08852_ (.A(_00950_),
    .B(_00951_),
    .Y(_00952_));
 sky130_fd_sc_hd__xor2_1 _08853_ (.A(_00949_),
    .B(_00952_),
    .X(_00953_));
 sky130_fd_sc_hd__nand2_1 _08854_ (.A(_00773_),
    .B(_00953_),
    .Y(_00954_));
 sky130_fd_sc_hd__or2_1 _08855_ (.A(_00773_),
    .B(_00953_),
    .X(_00955_));
 sky130_fd_sc_hd__nand2_1 _08856_ (.A(_00954_),
    .B(_00955_),
    .Y(_00957_));
 sky130_fd_sc_hd__and4_1 _08857_ (.A(_00431_),
    .B(_04169_),
    .C(net47),
    .D(net48),
    .X(_00958_));
 sky130_fd_sc_hd__clkbuf_4 _08858_ (.A(net48),
    .X(_00959_));
 sky130_fd_sc_hd__a22o_1 _08859_ (.A1(_03587_),
    .A2(net47),
    .B1(_00959_),
    .B2(_03576_),
    .X(_00960_));
 sky130_fd_sc_hd__or2b_1 _08860_ (.A(_00958_),
    .B_N(_00960_),
    .X(_00961_));
 sky130_fd_sc_hd__nand2_1 _08861_ (.A(_01372_),
    .B(net46),
    .Y(_00962_));
 sky130_fd_sc_hd__xnor2_1 _08862_ (.A(_00961_),
    .B(_00962_),
    .Y(_00963_));
 sky130_fd_sc_hd__a31o_1 _08863_ (.A1(_01284_),
    .A2(net45),
    .A3(_00793_),
    .B1(_00791_),
    .X(_00964_));
 sky130_fd_sc_hd__and2_1 _08864_ (.A(_01230_),
    .B(net45),
    .X(_00965_));
 sky130_fd_sc_hd__xnor2_1 _08865_ (.A(_00964_),
    .B(_00965_),
    .Y(_00966_));
 sky130_fd_sc_hd__xor2_1 _08866_ (.A(_00963_),
    .B(_00966_),
    .X(_00968_));
 sky130_fd_sc_hd__nand2_1 _08867_ (.A(_00797_),
    .B(_00968_),
    .Y(_00969_));
 sky130_fd_sc_hd__or2_1 _08868_ (.A(_00797_),
    .B(_00968_),
    .X(_00970_));
 sky130_fd_sc_hd__nand2_1 _08869_ (.A(_00969_),
    .B(_00970_),
    .Y(_00971_));
 sky130_fd_sc_hd__nand2_1 _08870_ (.A(_00776_),
    .B(_00786_),
    .Y(_00972_));
 sky130_fd_sc_hd__nand2_1 _08871_ (.A(_00787_),
    .B(_00788_),
    .Y(_00973_));
 sky130_fd_sc_hd__and3_1 _08872_ (.A(_00615_),
    .B(_00972_),
    .C(_00973_),
    .X(_00974_));
 sky130_fd_sc_hd__xor2_1 _08873_ (.A(_00971_),
    .B(_00974_),
    .X(_00975_));
 sky130_fd_sc_hd__xnor2_2 _08874_ (.A(_00957_),
    .B(_00975_),
    .Y(_00976_));
 sky130_fd_sc_hd__nor2_1 _08875_ (.A(_00789_),
    .B(_00799_),
    .Y(_00977_));
 sky130_fd_sc_hd__nand2_1 _08876_ (.A(_00789_),
    .B(_00799_),
    .Y(_00979_));
 sky130_fd_sc_hd__o21ai_1 _08877_ (.A1(_00775_),
    .A2(_00977_),
    .B1(_00979_),
    .Y(_00980_));
 sky130_fd_sc_hd__xnor2_2 _08878_ (.A(_00976_),
    .B(_00980_),
    .Y(_00981_));
 sky130_fd_sc_hd__and2b_1 _08879_ (.A_N(_00766_),
    .B(_00801_),
    .X(_00982_));
 sky130_fd_sc_hd__a21o_1 _08880_ (.A1(_00629_),
    .A2(_00802_),
    .B1(_00982_),
    .X(_00983_));
 sky130_fd_sc_hd__xnor2_2 _08881_ (.A(_00981_),
    .B(_00983_),
    .Y(_00984_));
 sky130_fd_sc_hd__nor2_1 _08882_ (.A(_00710_),
    .B(_00877_),
    .Y(_00985_));
 sky130_fd_sc_hd__and2_1 _08883_ (.A(_00713_),
    .B(_00985_),
    .X(_00986_));
 sky130_fd_sc_hd__nand2_1 _08884_ (.A(_00874_),
    .B(_00876_),
    .Y(_00987_));
 sky130_fd_sc_hd__nor2_1 _08885_ (.A(_00874_),
    .B(_00876_),
    .Y(_00988_));
 sky130_fd_sc_hd__a21oi_1 _08886_ (.A1(_00881_),
    .A2(_00987_),
    .B1(_00988_),
    .Y(_00990_));
 sky130_fd_sc_hd__a311o_4 _08887_ (.A1(_00251_),
    .A2(_00712_),
    .A3(_00985_),
    .B1(_00986_),
    .C1(_00990_),
    .X(_00991_));
 sky130_fd_sc_hd__or2b_1 _08888_ (.A(_00806_),
    .B_N(_00837_),
    .X(_00992_));
 sky130_fd_sc_hd__and4_1 _08889_ (.A(_06965_),
    .B(_06966_),
    .C(_04906_),
    .D(_04928_),
    .X(_00993_));
 sky130_fd_sc_hd__a22o_1 _08890_ (.A1(_06966_),
    .A2(_04906_),
    .B1(_04928_),
    .B2(_06965_),
    .X(_00994_));
 sky130_fd_sc_hd__and2b_1 _08891_ (.A_N(_00993_),
    .B(_00994_),
    .X(_00995_));
 sky130_fd_sc_hd__nand2_1 _08892_ (.A(_03543_),
    .B(_00144_),
    .Y(_00996_));
 sky130_fd_sc_hd__xnor2_1 _08893_ (.A(_00995_),
    .B(_00996_),
    .Y(_00997_));
 sky130_fd_sc_hd__o211ai_2 _08894_ (.A1(_00807_),
    .A2(_00809_),
    .B1(_00508_),
    .C1(_00298_),
    .Y(_00998_));
 sky130_fd_sc_hd__a211o_1 _08895_ (.A1(_00508_),
    .A2(_00158_),
    .B1(_00807_),
    .C1(_00809_),
    .X(_00999_));
 sky130_fd_sc_hd__and2_1 _08896_ (.A(_00998_),
    .B(_00999_),
    .X(_01001_));
 sky130_fd_sc_hd__nand2_1 _08897_ (.A(_00997_),
    .B(_01001_),
    .Y(_01002_));
 sky130_fd_sc_hd__or2_1 _08898_ (.A(_00997_),
    .B(_01001_),
    .X(_01003_));
 sky130_fd_sc_hd__nand2_1 _08899_ (.A(_01002_),
    .B(_01003_),
    .Y(_01004_));
 sky130_fd_sc_hd__nor2_1 _08900_ (.A(_00813_),
    .B(_01004_),
    .Y(_01005_));
 sky130_fd_sc_hd__and2_1 _08901_ (.A(_00813_),
    .B(_01004_),
    .X(_01006_));
 sky130_fd_sc_hd__or2_1 _08902_ (.A(_01005_),
    .B(_01006_),
    .X(_01007_));
 sky130_fd_sc_hd__and4_1 _08903_ (.A(_00377_),
    .B(_02993_),
    .C(_00112_),
    .D(_00268_),
    .X(_01008_));
 sky130_fd_sc_hd__a22oi_1 _08904_ (.A1(_00388_),
    .A2(_00112_),
    .B1(_00114_),
    .B2(_03004_),
    .Y(_01009_));
 sky130_fd_sc_hd__and4bb_1 _08905_ (.A_N(_01008_),
    .B_N(_01009_),
    .C(_06765_),
    .D(_00095_),
    .X(_01010_));
 sky130_fd_sc_hd__o2bb2a_1 _08906_ (.A1_N(_00003_),
    .A2_N(_00095_),
    .B1(_01008_),
    .B2(_01009_),
    .X(_01012_));
 sky130_fd_sc_hd__or2_1 _08907_ (.A(_01010_),
    .B(_01012_),
    .X(_01013_));
 sky130_fd_sc_hd__a32o_1 _08908_ (.A1(_06775_),
    .A2(_00095_),
    .A3(_00826_),
    .B1(_00656_),
    .B2(_00258_),
    .X(_01014_));
 sky130_fd_sc_hd__nand2_1 _08909_ (.A(_06775_),
    .B(_00151_),
    .Y(_01015_));
 sky130_fd_sc_hd__xnor2_1 _08910_ (.A(_01014_),
    .B(_01015_),
    .Y(_01016_));
 sky130_fd_sc_hd__xnor2_1 _08911_ (.A(_01013_),
    .B(_01016_),
    .Y(_01017_));
 sky130_fd_sc_hd__nand2_1 _08912_ (.A(_00830_),
    .B(_01017_),
    .Y(_01018_));
 sky130_fd_sc_hd__or2_1 _08913_ (.A(_00830_),
    .B(_01017_),
    .X(_01019_));
 sky130_fd_sc_hd__nand2_1 _08914_ (.A(_01018_),
    .B(_01019_),
    .Y(_01020_));
 sky130_fd_sc_hd__and2_1 _08915_ (.A(_00822_),
    .B(_00823_),
    .X(_01021_));
 sky130_fd_sc_hd__a211oi_2 _08916_ (.A1(_00817_),
    .A2(_00821_),
    .B1(_01021_),
    .C1(_00645_),
    .Y(_01023_));
 sky130_fd_sc_hd__xor2_1 _08917_ (.A(_01020_),
    .B(_01023_),
    .X(_01024_));
 sky130_fd_sc_hd__xnor2_1 _08918_ (.A(_01007_),
    .B(_01024_),
    .Y(_01025_));
 sky130_fd_sc_hd__nand2_1 _08919_ (.A(_00816_),
    .B(_00834_),
    .Y(_01026_));
 sky130_fd_sc_hd__and3_1 _08920_ (.A(_00833_),
    .B(_01025_),
    .C(_01026_),
    .X(_01027_));
 sky130_fd_sc_hd__a21oi_1 _08921_ (.A1(_00833_),
    .A2(_01026_),
    .B1(_01025_),
    .Y(_01028_));
 sky130_fd_sc_hd__or2_1 _08922_ (.A(_01027_),
    .B(_01028_),
    .X(_01029_));
 sky130_fd_sc_hd__a21oi_1 _08923_ (.A1(_00992_),
    .A2(_00839_),
    .B1(_01029_),
    .Y(_01030_));
 sky130_fd_sc_hd__and3_1 _08924_ (.A(_00992_),
    .B(_00839_),
    .C(_01029_),
    .X(_01031_));
 sky130_fd_sc_hd__or2_2 _08925_ (.A(_01030_),
    .B(_01031_),
    .X(_01032_));
 sky130_fd_sc_hd__and2_1 _08926_ (.A(_00857_),
    .B(_00871_),
    .X(_01034_));
 sky130_fd_sc_hd__or3_1 _08927_ (.A(_00673_),
    .B(_00848_),
    .C(_00852_),
    .X(_01035_));
 sky130_fd_sc_hd__a21oi_2 _08928_ (.A1(_00853_),
    .A2(_00856_),
    .B1(_01035_),
    .Y(_01036_));
 sky130_fd_sc_hd__inv_2 _08929_ (.A(_00866_),
    .Y(_01037_));
 sky130_fd_sc_hd__or3_1 _08930_ (.A(_00690_),
    .B(_00861_),
    .C(_00865_),
    .X(_01038_));
 sky130_fd_sc_hd__o21ba_2 _08931_ (.A1(_01037_),
    .A2(_00870_),
    .B1_N(_01038_),
    .X(_01039_));
 sky130_fd_sc_hd__xor2_2 _08932_ (.A(_01036_),
    .B(_01039_),
    .X(_01040_));
 sky130_fd_sc_hd__xor2_2 _08933_ (.A(_01034_),
    .B(_01040_),
    .X(_01041_));
 sky130_fd_sc_hd__xnor2_4 _08934_ (.A(_01032_),
    .B(_01041_),
    .Y(_01042_));
 sky130_fd_sc_hd__nor2_1 _08935_ (.A(_00842_),
    .B(_00872_),
    .Y(_01043_));
 sky130_fd_sc_hd__nand2_1 _08936_ (.A(_00842_),
    .B(_00872_),
    .Y(_01045_));
 sky130_fd_sc_hd__o21a_2 _08937_ (.A1(_00841_),
    .A2(_01043_),
    .B1(_01045_),
    .X(_01046_));
 sky130_fd_sc_hd__xnor2_4 _08938_ (.A(_01042_),
    .B(_01046_),
    .Y(_01047_));
 sky130_fd_sc_hd__xor2_2 _08939_ (.A(_00991_),
    .B(_01047_),
    .X(_01048_));
 sky130_fd_sc_hd__xor2_2 _08940_ (.A(_00984_),
    .B(_01048_),
    .X(_01049_));
 sky130_fd_sc_hd__xnor2_4 _08941_ (.A(_00943_),
    .B(_01049_),
    .Y(_01050_));
 sky130_fd_sc_hd__a21o_1 _08942_ (.A1(_00765_),
    .A2(_00887_),
    .B1(_00886_),
    .X(_01051_));
 sky130_fd_sc_hd__inv_2 _08943_ (.A(_01051_),
    .Y(_01052_));
 sky130_fd_sc_hd__xnor2_4 _08944_ (.A(_01050_),
    .B(_01052_),
    .Y(_01053_));
 sky130_fd_sc_hd__xnor2_4 _08945_ (.A(_00899_),
    .B(_01053_),
    .Y(_01054_));
 sky130_fd_sc_hd__xor2_2 _08946_ (.A(_00898_),
    .B(_01054_),
    .X(net80));
 sky130_fd_sc_hd__and2_4 _08947_ (.A(_01050_),
    .B(_01052_),
    .X(_01056_));
 sky130_fd_sc_hd__and2_1 _08948_ (.A(_00410_),
    .B(_00380_),
    .X(_01057_));
 sky130_fd_sc_hd__buf_2 _08949_ (.A(net49),
    .X(_01058_));
 sky130_fd_sc_hd__clkbuf_4 _08950_ (.A(_01058_),
    .X(_01059_));
 sky130_fd_sc_hd__clkbuf_4 _08951_ (.A(_01059_),
    .X(_01060_));
 sky130_fd_sc_hd__clkbuf_4 _08952_ (.A(_01060_),
    .X(_01061_));
 sky130_fd_sc_hd__buf_4 _08953_ (.A(_01061_),
    .X(_01062_));
 sky130_fd_sc_hd__o211a_1 _08954_ (.A1(_00775_),
    .A2(_00977_),
    .B1(_00976_),
    .C1(_00979_),
    .X(_01063_));
 sky130_fd_sc_hd__a21o_1 _08955_ (.A1(_00981_),
    .A2(_00983_),
    .B1(_01063_),
    .X(_01064_));
 sky130_fd_sc_hd__buf_4 _08956_ (.A(_00460_),
    .X(_01066_));
 sky130_fd_sc_hd__nand2_1 _08957_ (.A(_02467_),
    .B(_01066_),
    .Y(_01067_));
 sky130_fd_sc_hd__and2_1 _08958_ (.A(_00971_),
    .B(_00974_),
    .X(_01068_));
 sky130_fd_sc_hd__o21a_1 _08959_ (.A1(_00971_),
    .A2(_00974_),
    .B1(_00957_),
    .X(_01069_));
 sky130_fd_sc_hd__nand2_1 _08960_ (.A(_00964_),
    .B(_00965_),
    .Y(_01070_));
 sky130_fd_sc_hd__o21a_1 _08961_ (.A1(_00963_),
    .A2(_00966_),
    .B1(_01070_),
    .X(_01071_));
 sky130_fd_sc_hd__a31o_1 _08962_ (.A1(_04081_),
    .A2(_00604_),
    .A3(_00960_),
    .B1(_00958_),
    .X(_01072_));
 sky130_fd_sc_hd__and4_1 _08963_ (.A(_04169_),
    .B(_01076_),
    .C(net47),
    .D(net48),
    .X(_01073_));
 sky130_fd_sc_hd__a22o_1 _08964_ (.A1(_01076_),
    .A2(net47),
    .B1(_00959_),
    .B2(_03587_),
    .X(_01074_));
 sky130_fd_sc_hd__and2b_1 _08965_ (.A_N(_01073_),
    .B(_01074_),
    .X(_01075_));
 sky130_fd_sc_hd__nand2_1 _08966_ (.A(_04268_),
    .B(net46),
    .Y(_01077_));
 sky130_fd_sc_hd__xnor2_2 _08967_ (.A(_01075_),
    .B(_01077_),
    .Y(_01078_));
 sky130_fd_sc_hd__xor2_1 _08968_ (.A(_01072_),
    .B(_01078_),
    .X(_01079_));
 sky130_fd_sc_hd__xor2_1 _08969_ (.A(_01071_),
    .B(_01079_),
    .X(_01080_));
 sky130_fd_sc_hd__nor2_1 _08970_ (.A(_00969_),
    .B(_01080_),
    .Y(_01081_));
 sky130_fd_sc_hd__and2_1 _08971_ (.A(_00969_),
    .B(_01080_),
    .X(_01082_));
 sky130_fd_sc_hd__nor2_1 _08972_ (.A(_01081_),
    .B(_01082_),
    .Y(_01083_));
 sky130_fd_sc_hd__nand2_1 _08973_ (.A(_00950_),
    .B(_00951_),
    .Y(_01084_));
 sky130_fd_sc_hd__o21a_1 _08974_ (.A1(_00949_),
    .A2(_00952_),
    .B1(_01084_),
    .X(_01085_));
 sky130_fd_sc_hd__a31o_1 _08975_ (.A1(_05577_),
    .A2(_00373_),
    .A3(_00946_),
    .B1(_00944_),
    .X(_01086_));
 sky130_fd_sc_hd__and4_1 _08976_ (.A(_00639_),
    .B(net29),
    .C(_04180_),
    .D(_04191_),
    .X(_01088_));
 sky130_fd_sc_hd__a22o_1 _08977_ (.A1(_00541_),
    .A2(_04103_),
    .B1(_04191_),
    .B2(_00639_),
    .X(_01089_));
 sky130_fd_sc_hd__and2b_1 _08978_ (.A_N(_01088_),
    .B(_01089_),
    .X(_01090_));
 sky130_fd_sc_hd__nand2_1 _08979_ (.A(_03268_),
    .B(_04026_),
    .Y(_01091_));
 sky130_fd_sc_hd__xnor2_1 _08980_ (.A(_01090_),
    .B(_01091_),
    .Y(_01092_));
 sky130_fd_sc_hd__xor2_1 _08981_ (.A(_01086_),
    .B(_01092_),
    .X(_01093_));
 sky130_fd_sc_hd__xor2_1 _08982_ (.A(_01085_),
    .B(_01093_),
    .X(_01094_));
 sky130_fd_sc_hd__nor2_1 _08983_ (.A(_00954_),
    .B(_01094_),
    .Y(_01095_));
 sky130_fd_sc_hd__and2_1 _08984_ (.A(_00954_),
    .B(_01094_),
    .X(_01096_));
 sky130_fd_sc_hd__nor2_1 _08985_ (.A(_01095_),
    .B(_01096_),
    .Y(_01097_));
 sky130_fd_sc_hd__nand2_1 _08986_ (.A(_01083_),
    .B(_01097_),
    .Y(_01099_));
 sky130_fd_sc_hd__or2_1 _08987_ (.A(_01083_),
    .B(_01097_),
    .X(_01100_));
 sky130_fd_sc_hd__nand2_1 _08988_ (.A(_01099_),
    .B(_01100_),
    .Y(_01101_));
 sky130_fd_sc_hd__o21a_1 _08989_ (.A1(_01068_),
    .A2(_01069_),
    .B1(_01101_),
    .X(_01102_));
 sky130_fd_sc_hd__or3_1 _08990_ (.A(_01068_),
    .B(_01101_),
    .C(_01069_),
    .X(_01103_));
 sky130_fd_sc_hd__and2b_1 _08991_ (.A_N(_01102_),
    .B(_01103_),
    .X(_01104_));
 sky130_fd_sc_hd__xnor2_2 _08992_ (.A(_01067_),
    .B(_01104_),
    .Y(_01105_));
 sky130_fd_sc_hd__xor2_1 _08993_ (.A(_01064_),
    .B(_01105_),
    .X(_01106_));
 sky130_fd_sc_hd__and3_1 _08994_ (.A(_00464_),
    .B(_01062_),
    .C(_01106_),
    .X(_01107_));
 sky130_fd_sc_hd__clkbuf_8 _08995_ (.A(_01062_),
    .X(_01108_));
 sky130_fd_sc_hd__a21o_1 _08996_ (.A1(_00464_),
    .A2(_01108_),
    .B1(_01106_),
    .X(_01110_));
 sky130_fd_sc_hd__or2b_1 _08997_ (.A(_01107_),
    .B_N(_01110_),
    .X(_01111_));
 sky130_fd_sc_hd__xnor2_2 _08998_ (.A(_01057_),
    .B(_01111_),
    .Y(_01112_));
 sky130_fd_sc_hd__or2_1 _08999_ (.A(_01034_),
    .B(_01040_),
    .X(_01113_));
 sky130_fd_sc_hd__a21bo_1 _09000_ (.A1(_01034_),
    .A2(_01040_),
    .B1_N(_01032_),
    .X(_01114_));
 sky130_fd_sc_hd__nor2_1 _09001_ (.A(_01036_),
    .B(_01039_),
    .Y(_01115_));
 sky130_fd_sc_hd__nor2_1 _09002_ (.A(_01027_),
    .B(_01030_),
    .Y(_01116_));
 sky130_fd_sc_hd__and2_1 _09003_ (.A(_01020_),
    .B(_01023_),
    .X(_01117_));
 sky130_fd_sc_hd__o21a_1 _09004_ (.A1(_01020_),
    .A2(_01023_),
    .B1(_01007_),
    .X(_01118_));
 sky130_fd_sc_hd__and3_1 _09005_ (.A(_06885_),
    .B(_00294_),
    .C(_01014_),
    .X(_01119_));
 sky130_fd_sc_hd__and2b_1 _09006_ (.A_N(_01013_),
    .B(_01016_),
    .X(_01121_));
 sky130_fd_sc_hd__nor2_1 _09007_ (.A(_01008_),
    .B(_01010_),
    .Y(_01122_));
 sky130_fd_sc_hd__a22oi_2 _09008_ (.A1(_03004_),
    .A2(_00113_),
    .B1(_00114_),
    .B2(_00095_),
    .Y(_01123_));
 sky130_fd_sc_hd__and4_1 _09009_ (.A(_03004_),
    .B(_00113_),
    .C(_00114_),
    .D(_00094_),
    .X(_01124_));
 sky130_fd_sc_hd__nor2_1 _09010_ (.A(_01123_),
    .B(_01124_),
    .Y(_01125_));
 sky130_fd_sc_hd__nand2_1 _09011_ (.A(_00003_),
    .B(_00151_),
    .Y(_01126_));
 sky130_fd_sc_hd__xnor2_1 _09012_ (.A(_01125_),
    .B(_01126_),
    .Y(_01127_));
 sky130_fd_sc_hd__xnor2_1 _09013_ (.A(_01122_),
    .B(_01127_),
    .Y(_01128_));
 sky130_fd_sc_hd__o21ai_1 _09014_ (.A1(_01119_),
    .A2(_01121_),
    .B1(_01128_),
    .Y(_01129_));
 sky130_fd_sc_hd__or3_1 _09015_ (.A(_01119_),
    .B(_01121_),
    .C(_01128_),
    .X(_01130_));
 sky130_fd_sc_hd__nand2_1 _09016_ (.A(_01129_),
    .B(_01130_),
    .Y(_01132_));
 sky130_fd_sc_hd__xor2_1 _09017_ (.A(_01018_),
    .B(_01132_),
    .X(_01133_));
 sky130_fd_sc_hd__a31o_1 _09018_ (.A1(_03543_),
    .A2(_00144_),
    .A3(_00994_),
    .B1(_00993_),
    .X(_01134_));
 sky130_fd_sc_hd__nand2_1 _09019_ (.A(_06965_),
    .B(_04906_),
    .Y(_01135_));
 sky130_fd_sc_hd__nand2_1 _09020_ (.A(_06966_),
    .B(_00142_),
    .Y(_01136_));
 sky130_fd_sc_hd__and4_1 _09021_ (.A(_06964_),
    .B(_06966_),
    .C(_00142_),
    .D(_04895_),
    .X(_01137_));
 sky130_fd_sc_hd__a21oi_1 _09022_ (.A1(_01135_),
    .A2(_01136_),
    .B1(_01137_),
    .Y(_01138_));
 sky130_fd_sc_hd__a21oi_1 _09023_ (.A1(_03543_),
    .A2(_00298_),
    .B1(_01138_),
    .Y(_01139_));
 sky130_fd_sc_hd__and3_1 _09024_ (.A(_03543_),
    .B(_00298_),
    .C(_01138_),
    .X(_01140_));
 sky130_fd_sc_hd__nor2_1 _09025_ (.A(_01139_),
    .B(_01140_),
    .Y(_01141_));
 sky130_fd_sc_hd__xnor2_1 _09026_ (.A(_01134_),
    .B(_01141_),
    .Y(_01143_));
 sky130_fd_sc_hd__a21o_1 _09027_ (.A1(_00998_),
    .A2(_01002_),
    .B1(_01143_),
    .X(_01144_));
 sky130_fd_sc_hd__nand3_1 _09028_ (.A(_00998_),
    .B(_01002_),
    .C(_01143_),
    .Y(_01145_));
 sky130_fd_sc_hd__and2_1 _09029_ (.A(_01144_),
    .B(_01145_),
    .X(_01146_));
 sky130_fd_sc_hd__xnor2_1 _09030_ (.A(_01005_),
    .B(_01146_),
    .Y(_01147_));
 sky130_fd_sc_hd__inv_2 _09031_ (.A(_01147_),
    .Y(_01148_));
 sky130_fd_sc_hd__nand2_1 _09032_ (.A(_01133_),
    .B(_01148_),
    .Y(_01149_));
 sky130_fd_sc_hd__or2_1 _09033_ (.A(_01133_),
    .B(_01148_),
    .X(_01150_));
 sky130_fd_sc_hd__nand2_1 _09034_ (.A(_01149_),
    .B(_01150_),
    .Y(_01151_));
 sky130_fd_sc_hd__o21a_1 _09035_ (.A1(_01117_),
    .A2(_01118_),
    .B1(_01151_),
    .X(_01152_));
 sky130_fd_sc_hd__nor3_1 _09036_ (.A(_01117_),
    .B(_01151_),
    .C(_01118_),
    .Y(_01154_));
 sky130_fd_sc_hd__buf_4 _09037_ (.A(_00544_),
    .X(_01155_));
 sky130_fd_sc_hd__clkbuf_4 _09038_ (.A(_00526_),
    .X(_01156_));
 sky130_fd_sc_hd__o211ai_1 _09039_ (.A1(_01152_),
    .A2(_01154_),
    .B1(_01155_),
    .C1(_01156_),
    .Y(_01157_));
 sky130_fd_sc_hd__a211o_1 _09040_ (.A1(_01155_),
    .A2(_01156_),
    .B1(_01152_),
    .C1(_01154_),
    .X(_01158_));
 sky130_fd_sc_hd__nand2_2 _09041_ (.A(_01157_),
    .B(_01158_),
    .Y(_01159_));
 sky130_fd_sc_hd__xnor2_2 _09042_ (.A(_01116_),
    .B(_01159_),
    .Y(_01160_));
 sky130_fd_sc_hd__xor2_1 _09043_ (.A(_01115_),
    .B(_01160_),
    .X(_01161_));
 sky130_fd_sc_hd__a21o_1 _09044_ (.A1(_01113_),
    .A2(_01114_),
    .B1(_01161_),
    .X(_01162_));
 sky130_fd_sc_hd__and3_1 _09045_ (.A(_01113_),
    .B(_01161_),
    .C(_01114_),
    .X(_01163_));
 sky130_fd_sc_hd__inv_2 _09046_ (.A(_01163_),
    .Y(_01165_));
 sky130_fd_sc_hd__and2_1 _09047_ (.A(_01162_),
    .B(_01165_),
    .X(_01166_));
 sky130_fd_sc_hd__nor3_2 _09048_ (.A(_00877_),
    .B(_00878_),
    .C(_01047_),
    .Y(_01167_));
 sky130_fd_sc_hd__nand2_1 _09049_ (.A(_01042_),
    .B(_01046_),
    .Y(_01168_));
 sky130_fd_sc_hd__or2_1 _09050_ (.A(_01042_),
    .B(_01046_),
    .X(_01169_));
 sky130_fd_sc_hd__a21bo_1 _09051_ (.A1(_00987_),
    .A2(_01168_),
    .B1_N(_01169_),
    .X(_01170_));
 sky130_fd_sc_hd__a2111o_1 _09052_ (.A1(_00711_),
    .A2(_00881_),
    .B1(_00882_),
    .C1(_00877_),
    .D1(_01047_),
    .X(_01171_));
 sky130_fd_sc_hd__nand2_1 _09053_ (.A(_01170_),
    .B(_01171_),
    .Y(_01172_));
 sky130_fd_sc_hd__a21o_1 _09054_ (.A1(_00557_),
    .A2(_01167_),
    .B1(_01172_),
    .X(_01173_));
 sky130_fd_sc_hd__xor2_2 _09055_ (.A(_01166_),
    .B(_01173_),
    .X(_01174_));
 sky130_fd_sc_hd__xnor2_2 _09056_ (.A(_01112_),
    .B(_01174_),
    .Y(_01176_));
 sky130_fd_sc_hd__clkbuf_4 _09057_ (.A(net17),
    .X(_01177_));
 sky130_fd_sc_hd__clkbuf_4 _09058_ (.A(_01177_),
    .X(_01178_));
 sky130_fd_sc_hd__buf_4 _09059_ (.A(_01178_),
    .X(_01179_));
 sky130_fd_sc_hd__buf_4 _09060_ (.A(_01179_),
    .X(_01180_));
 sky130_fd_sc_hd__clkbuf_4 _09061_ (.A(_01180_),
    .X(_01181_));
 sky130_fd_sc_hd__buf_4 _09062_ (.A(_01181_),
    .X(_01182_));
 sky130_fd_sc_hd__buf_4 _09063_ (.A(_01182_),
    .X(_01183_));
 sky130_fd_sc_hd__nand2_2 _09064_ (.A(_00344_),
    .B(_01183_),
    .Y(_01184_));
 sky130_fd_sc_hd__o211a_1 _09065_ (.A1(_00740_),
    .A2(_00937_),
    .B1(_00936_),
    .C1(_00938_),
    .X(_01185_));
 sky130_fd_sc_hd__a21o_1 _09066_ (.A1(_00940_),
    .A2(_00942_),
    .B1(_01185_),
    .X(_01187_));
 sky130_fd_sc_hd__buf_4 _09067_ (.A(_00416_),
    .X(_01188_));
 sky130_fd_sc_hd__nand2_1 _09068_ (.A(_02456_),
    .B(_01188_),
    .Y(_01189_));
 sky130_fd_sc_hd__nand2_1 _09069_ (.A(_00913_),
    .B(_00933_),
    .Y(_01190_));
 sky130_fd_sc_hd__nand2_1 _09070_ (.A(_00925_),
    .B(_00926_),
    .Y(_01191_));
 sky130_fd_sc_hd__a21bo_1 _09071_ (.A1(_00924_),
    .A2(_00927_),
    .B1_N(_01191_),
    .X(_01192_));
 sky130_fd_sc_hd__a31o_1 _09072_ (.A1(_01996_),
    .A2(_03894_),
    .A3(_00920_),
    .B1(_00919_),
    .X(_01193_));
 sky130_fd_sc_hd__and4_1 _09073_ (.A(_05445_),
    .B(_05731_),
    .C(_03718_),
    .D(net10),
    .X(_01194_));
 sky130_fd_sc_hd__a22oi_1 _09074_ (.A1(_05445_),
    .A2(_00423_),
    .B1(net10),
    .B2(_05731_),
    .Y(_01195_));
 sky130_fd_sc_hd__and4bb_1 _09075_ (.A_N(_01194_),
    .B_N(_01195_),
    .C(_01996_),
    .D(net11),
    .X(_01196_));
 sky130_fd_sc_hd__o2bb2a_1 _09076_ (.A1_N(_01996_),
    .A2_N(net11),
    .B1(_01194_),
    .B2(_01195_),
    .X(_01198_));
 sky130_fd_sc_hd__nor2_1 _09077_ (.A(_01196_),
    .B(_01198_),
    .Y(_01199_));
 sky130_fd_sc_hd__xor2_1 _09078_ (.A(_01193_),
    .B(_01199_),
    .X(_01200_));
 sky130_fd_sc_hd__xor2_1 _09079_ (.A(_01192_),
    .B(_01200_),
    .X(_01201_));
 sky130_fd_sc_hd__nand2_1 _09080_ (.A(_00929_),
    .B(_01201_),
    .Y(_01202_));
 sky130_fd_sc_hd__or2_1 _09081_ (.A(_00929_),
    .B(_01201_),
    .X(_01203_));
 sky130_fd_sc_hd__nand2_1 _09082_ (.A(_01202_),
    .B(_01203_),
    .Y(_01204_));
 sky130_fd_sc_hd__nand2_1 _09083_ (.A(_00906_),
    .B(_00907_),
    .Y(_01205_));
 sky130_fd_sc_hd__a21bo_1 _09084_ (.A1(_00905_),
    .A2(_00908_),
    .B1_N(_01205_),
    .X(_01206_));
 sky130_fd_sc_hd__a31o_1 _09085_ (.A1(_02127_),
    .A2(_00734_),
    .A3(_00902_),
    .B1(_00900_),
    .X(_01207_));
 sky130_fd_sc_hd__and4_1 _09086_ (.A(_03850_),
    .B(_01394_),
    .C(_00730_),
    .D(net15),
    .X(_01209_));
 sky130_fd_sc_hd__a22oi_1 _09087_ (.A1(_03850_),
    .A2(_00730_),
    .B1(net15),
    .B2(_01306_),
    .Y(_01210_));
 sky130_fd_sc_hd__clkbuf_4 _09088_ (.A(net16),
    .X(_01211_));
 sky130_fd_sc_hd__and4bb_1 _09089_ (.A_N(_01209_),
    .B_N(_01210_),
    .C(_01744_),
    .D(_01211_),
    .X(_01212_));
 sky130_fd_sc_hd__o2bb2a_1 _09090_ (.A1_N(_01744_),
    .A2_N(_01211_),
    .B1(_01209_),
    .B2(_01210_),
    .X(_01213_));
 sky130_fd_sc_hd__nor2_1 _09091_ (.A(_01212_),
    .B(_01213_),
    .Y(_01214_));
 sky130_fd_sc_hd__xor2_1 _09092_ (.A(_01207_),
    .B(_01214_),
    .X(_01215_));
 sky130_fd_sc_hd__xor2_1 _09093_ (.A(_01206_),
    .B(_01215_),
    .X(_01216_));
 sky130_fd_sc_hd__nand2_1 _09094_ (.A(_00910_),
    .B(_01216_),
    .Y(_01217_));
 sky130_fd_sc_hd__or2_1 _09095_ (.A(_00910_),
    .B(_01216_),
    .X(_01218_));
 sky130_fd_sc_hd__nand2_1 _09096_ (.A(_01217_),
    .B(_01218_),
    .Y(_01220_));
 sky130_fd_sc_hd__nor2_1 _09097_ (.A(_01204_),
    .B(_01220_),
    .Y(_01221_));
 sky130_fd_sc_hd__and2_1 _09098_ (.A(_01204_),
    .B(_01220_),
    .X(_01222_));
 sky130_fd_sc_hd__nor2_1 _09099_ (.A(_01221_),
    .B(_01222_),
    .Y(_01223_));
 sky130_fd_sc_hd__a21oi_1 _09100_ (.A1(_00932_),
    .A2(_01190_),
    .B1(_01223_),
    .Y(_01224_));
 sky130_fd_sc_hd__nand3_1 _09101_ (.A(_00932_),
    .B(_01223_),
    .C(_01190_),
    .Y(_01225_));
 sky130_fd_sc_hd__or2b_1 _09102_ (.A(_01224_),
    .B_N(_01225_),
    .X(_01226_));
 sky130_fd_sc_hd__xor2_2 _09103_ (.A(_01189_),
    .B(_01226_),
    .X(_01227_));
 sky130_fd_sc_hd__xor2_1 _09104_ (.A(_01187_),
    .B(_01227_),
    .X(_01228_));
 sky130_fd_sc_hd__and3_1 _09105_ (.A(_00530_),
    .B(_00391_),
    .C(_01228_),
    .X(_01229_));
 sky130_fd_sc_hd__a21o_1 _09106_ (.A1(_00530_),
    .A2(_00391_),
    .B1(_01228_),
    .X(_01231_));
 sky130_fd_sc_hd__or2b_2 _09107_ (.A(_01229_),
    .B_N(_01231_),
    .X(_01232_));
 sky130_fd_sc_hd__xnor2_4 _09108_ (.A(_01184_),
    .B(_01232_),
    .Y(_01233_));
 sky130_fd_sc_hd__xnor2_4 _09109_ (.A(_01176_),
    .B(_01233_),
    .Y(_01234_));
 sky130_fd_sc_hd__or2_1 _09110_ (.A(_00984_),
    .B(_01048_),
    .X(_01235_));
 sky130_fd_sc_hd__and2_1 _09111_ (.A(_00984_),
    .B(_01048_),
    .X(_01236_));
 sky130_fd_sc_hd__a21oi_4 _09112_ (.A1(_00943_),
    .A2(_01235_),
    .B1(_01236_),
    .Y(_01237_));
 sky130_fd_sc_hd__xnor2_4 _09113_ (.A(_01234_),
    .B(_01237_),
    .Y(_01238_));
 sky130_fd_sc_hd__xnor2_4 _09114_ (.A(_01056_),
    .B(_01238_),
    .Y(_01239_));
 sky130_fd_sc_hd__a21boi_1 _09115_ (.A1(_00727_),
    .A2(_00893_),
    .B1_N(_00899_),
    .Y(_01240_));
 sky130_fd_sc_hd__o32ai_2 _09116_ (.A1(_00894_),
    .A2(_00896_),
    .A3(_01054_),
    .B1(_01240_),
    .B2(_01053_),
    .Y(_01242_));
 sky130_fd_sc_hd__xnor2_4 _09117_ (.A(_01239_),
    .B(net131),
    .Y(net81));
 sky130_fd_sc_hd__nor2b_4 _09118_ (.A(_01234_),
    .B_N(_01237_),
    .Y(_01243_));
 sky130_fd_sc_hd__a21o_1 _09119_ (.A1(_00344_),
    .A2(_01182_),
    .B1(_01229_),
    .X(_01244_));
 sky130_fd_sc_hd__nand2_1 _09120_ (.A(_01231_),
    .B(_01244_),
    .Y(_01245_));
 sky130_fd_sc_hd__buf_2 _09121_ (.A(net18),
    .X(_01246_));
 sky130_fd_sc_hd__buf_2 _09122_ (.A(_01246_),
    .X(_01247_));
 sky130_fd_sc_hd__buf_2 _09123_ (.A(_01247_),
    .X(_01248_));
 sky130_fd_sc_hd__buf_4 _09124_ (.A(_01248_),
    .X(_01249_));
 sky130_fd_sc_hd__clkbuf_4 _09125_ (.A(_01249_),
    .X(_01250_));
 sky130_fd_sc_hd__buf_4 _09126_ (.A(_01250_),
    .X(_01252_));
 sky130_fd_sc_hd__a22o_1 _09127_ (.A1(_02138_),
    .A2(_01182_),
    .B1(_01252_),
    .B2(_00344_),
    .X(_01253_));
 sky130_fd_sc_hd__clkbuf_4 _09128_ (.A(_01247_),
    .X(_01254_));
 sky130_fd_sc_hd__nand4_4 _09129_ (.A(_02138_),
    .B(_00322_),
    .C(_01179_),
    .D(_01254_),
    .Y(_01255_));
 sky130_fd_sc_hd__and2_1 _09130_ (.A(_01253_),
    .B(_01255_),
    .X(_01256_));
 sky130_fd_sc_hd__nand2_1 _09131_ (.A(_01192_),
    .B(_01200_),
    .Y(_01257_));
 sky130_fd_sc_hd__nand2_1 _09132_ (.A(_01193_),
    .B(_01199_),
    .Y(_01258_));
 sky130_fd_sc_hd__a22o_1 _09133_ (.A1(_05456_),
    .A2(_03773_),
    .B1(_03938_),
    .B2(_05467_),
    .X(_01259_));
 sky130_fd_sc_hd__clkbuf_4 _09134_ (.A(_03938_),
    .X(_01260_));
 sky130_fd_sc_hd__nand4_2 _09135_ (.A(_05456_),
    .B(_05478_),
    .C(_03773_),
    .D(_01260_),
    .Y(_01261_));
 sky130_fd_sc_hd__o211a_1 _09136_ (.A1(_01194_),
    .A2(_01196_),
    .B1(_01259_),
    .C1(_01261_),
    .X(_01263_));
 sky130_fd_sc_hd__a211oi_1 _09137_ (.A1(_01259_),
    .A2(_01261_),
    .B1(_01194_),
    .C1(_01196_),
    .Y(_01264_));
 sky130_fd_sc_hd__nor2_1 _09138_ (.A(_01263_),
    .B(_01264_),
    .Y(_01265_));
 sky130_fd_sc_hd__xor2_1 _09139_ (.A(_01258_),
    .B(_01265_),
    .X(_01266_));
 sky130_fd_sc_hd__a21oi_1 _09140_ (.A1(_01257_),
    .A2(_01202_),
    .B1(_01266_),
    .Y(_01267_));
 sky130_fd_sc_hd__and3_1 _09141_ (.A(_01257_),
    .B(_01202_),
    .C(_01266_),
    .X(_01268_));
 sky130_fd_sc_hd__nor2_1 _09142_ (.A(_01267_),
    .B(_01268_),
    .Y(_01269_));
 sky130_fd_sc_hd__nand2_1 _09143_ (.A(_01206_),
    .B(_01215_),
    .Y(_01270_));
 sky130_fd_sc_hd__nand2_1 _09144_ (.A(_01207_),
    .B(_01214_),
    .Y(_01271_));
 sky130_fd_sc_hd__clkbuf_4 _09145_ (.A(net15),
    .X(_01272_));
 sky130_fd_sc_hd__a22o_1 _09146_ (.A1(_01295_),
    .A2(_01272_),
    .B1(_01211_),
    .B2(_01405_),
    .X(_01274_));
 sky130_fd_sc_hd__nand4_1 _09147_ (.A(_01361_),
    .B(_01405_),
    .C(_01272_),
    .D(_01211_),
    .Y(_01275_));
 sky130_fd_sc_hd__o211a_1 _09148_ (.A1(_01209_),
    .A2(_01212_),
    .B1(_01274_),
    .C1(_01275_),
    .X(_01276_));
 sky130_fd_sc_hd__a211oi_1 _09149_ (.A1(_01274_),
    .A2(_01275_),
    .B1(_01209_),
    .C1(_01212_),
    .Y(_01277_));
 sky130_fd_sc_hd__nor2_1 _09150_ (.A(_01276_),
    .B(_01277_),
    .Y(_01278_));
 sky130_fd_sc_hd__xor2_1 _09151_ (.A(_01271_),
    .B(_01278_),
    .X(_01279_));
 sky130_fd_sc_hd__a21oi_1 _09152_ (.A1(_01270_),
    .A2(_01217_),
    .B1(_01279_),
    .Y(_01280_));
 sky130_fd_sc_hd__and3_1 _09153_ (.A(_01270_),
    .B(_01217_),
    .C(_01279_),
    .X(_01281_));
 sky130_fd_sc_hd__nor2_1 _09154_ (.A(_01280_),
    .B(_01281_),
    .Y(_01282_));
 sky130_fd_sc_hd__xor2_1 _09155_ (.A(_01269_),
    .B(_01282_),
    .X(_01283_));
 sky130_fd_sc_hd__or2_1 _09156_ (.A(_01221_),
    .B(_01283_),
    .X(_01285_));
 sky130_fd_sc_hd__nand2_1 _09157_ (.A(_01221_),
    .B(_01283_),
    .Y(_01286_));
 sky130_fd_sc_hd__nand2_1 _09158_ (.A(_01285_),
    .B(_01286_),
    .Y(_01287_));
 sky130_fd_sc_hd__clkbuf_4 _09159_ (.A(_00575_),
    .X(_01288_));
 sky130_fd_sc_hd__buf_4 _09160_ (.A(_01288_),
    .X(_01289_));
 sky130_fd_sc_hd__a22o_1 _09161_ (.A1(_03070_),
    .A2(_01188_),
    .B1(_01289_),
    .B2(_02456_),
    .X(_01290_));
 sky130_fd_sc_hd__and4_1 _09162_ (.A(_03070_),
    .B(_02280_),
    .C(_00416_),
    .D(_01288_),
    .X(_01291_));
 sky130_fd_sc_hd__inv_2 _09163_ (.A(_01291_),
    .Y(_01292_));
 sky130_fd_sc_hd__and2_1 _09164_ (.A(_01290_),
    .B(_01292_),
    .X(_01293_));
 sky130_fd_sc_hd__xnor2_1 _09165_ (.A(_01287_),
    .B(_01293_),
    .Y(_01294_));
 sky130_fd_sc_hd__a21o_1 _09166_ (.A1(_01189_),
    .A2(_01225_),
    .B1(_01224_),
    .X(_01296_));
 sky130_fd_sc_hd__xnor2_1 _09167_ (.A(_01294_),
    .B(_01296_),
    .Y(_01297_));
 sky130_fd_sc_hd__and3_1 _09168_ (.A(_01187_),
    .B(_01227_),
    .C(_01297_),
    .X(_01298_));
 sky130_fd_sc_hd__a21oi_1 _09169_ (.A1(_01187_),
    .A2(_01227_),
    .B1(_01297_),
    .Y(_01299_));
 sky130_fd_sc_hd__nor2_1 _09170_ (.A(_01298_),
    .B(_01299_),
    .Y(_01300_));
 sky130_fd_sc_hd__a22o_1 _09171_ (.A1(_03554_),
    .A2(_00391_),
    .B1(_00393_),
    .B2(_00519_),
    .X(_01301_));
 sky130_fd_sc_hd__nand4_4 _09172_ (.A(_03521_),
    .B(_00486_),
    .C(_03707_),
    .D(_03740_),
    .Y(_01302_));
 sky130_fd_sc_hd__nand2_1 _09173_ (.A(_01301_),
    .B(_01302_),
    .Y(_01303_));
 sky130_fd_sc_hd__xnor2_1 _09174_ (.A(_01300_),
    .B(_01303_),
    .Y(_01304_));
 sky130_fd_sc_hd__xnor2_2 _09175_ (.A(_01256_),
    .B(_01304_),
    .Y(_01305_));
 sky130_fd_sc_hd__nor2_4 _09176_ (.A(_01245_),
    .B(_01305_),
    .Y(_01307_));
 sky130_fd_sc_hd__and2_1 _09177_ (.A(_01245_),
    .B(_01305_),
    .X(_01308_));
 sky130_fd_sc_hd__nor2_4 _09178_ (.A(_01307_),
    .B(_01308_),
    .Y(_01309_));
 sky130_fd_sc_hd__nand2_1 _09179_ (.A(_01115_),
    .B(_01160_),
    .Y(_01310_));
 sky130_fd_sc_hd__o21ai_2 _09180_ (.A1(_01027_),
    .A2(_01030_),
    .B1(_01159_),
    .Y(_01311_));
 sky130_fd_sc_hd__clkbuf_4 _09181_ (.A(_00654_),
    .X(_01312_));
 sky130_fd_sc_hd__a22o_1 _09182_ (.A1(_00544_),
    .A2(_00636_),
    .B1(_00526_),
    .B2(_01312_),
    .X(_01313_));
 sky130_fd_sc_hd__and4_1 _09183_ (.A(_01312_),
    .B(_00543_),
    .C(_00636_),
    .D(_00526_),
    .X(_01314_));
 sky130_fd_sc_hd__inv_2 _09184_ (.A(_01314_),
    .Y(_01315_));
 sky130_fd_sc_hd__and2_1 _09185_ (.A(_01313_),
    .B(_01315_),
    .X(_01316_));
 sky130_fd_sc_hd__or2b_1 _09186_ (.A(_01122_),
    .B_N(_01127_),
    .X(_01318_));
 sky130_fd_sc_hd__o21ba_1 _09187_ (.A1(_01123_),
    .A2(_01126_),
    .B1_N(_01124_),
    .X(_01319_));
 sky130_fd_sc_hd__a22o_1 _09188_ (.A1(_00257_),
    .A2(_00293_),
    .B1(_00294_),
    .B2(_00670_),
    .X(_01320_));
 sky130_fd_sc_hd__nand4_1 _09189_ (.A(_00257_),
    .B(_00670_),
    .C(_00819_),
    .D(_00818_),
    .Y(_01321_));
 sky130_fd_sc_hd__nand2_1 _09190_ (.A(_01320_),
    .B(_01321_),
    .Y(_01322_));
 sky130_fd_sc_hd__xor2_1 _09191_ (.A(_01319_),
    .B(_01322_),
    .X(_01323_));
 sky130_fd_sc_hd__xnor2_1 _09192_ (.A(_01318_),
    .B(_01323_),
    .Y(_01324_));
 sky130_fd_sc_hd__o21a_1 _09193_ (.A1(_01018_),
    .A2(_01132_),
    .B1(_01129_),
    .X(_01325_));
 sky130_fd_sc_hd__and2b_1 _09194_ (.A_N(_01324_),
    .B(_01325_),
    .X(_01326_));
 sky130_fd_sc_hd__and2b_1 _09195_ (.A_N(_01325_),
    .B(_01324_),
    .X(_01327_));
 sky130_fd_sc_hd__nor2_1 _09196_ (.A(_01326_),
    .B(_01327_),
    .Y(_01329_));
 sky130_fd_sc_hd__nand2_1 _09197_ (.A(_01005_),
    .B(_01146_),
    .Y(_01330_));
 sky130_fd_sc_hd__and2_1 _09198_ (.A(_01134_),
    .B(_01141_),
    .X(_01331_));
 sky130_fd_sc_hd__nor2_1 _09199_ (.A(_01137_),
    .B(_01140_),
    .Y(_01332_));
 sky130_fd_sc_hd__a22oi_1 _09200_ (.A1(_00262_),
    .A2(_00144_),
    .B1(_00298_),
    .B2(_00263_),
    .Y(_01333_));
 sky130_fd_sc_hd__and4_1 _09201_ (.A(_06965_),
    .B(_06966_),
    .C(_00143_),
    .D(_00158_),
    .X(_01334_));
 sky130_fd_sc_hd__or2_1 _09202_ (.A(_01333_),
    .B(_01334_),
    .X(_01335_));
 sky130_fd_sc_hd__xor2_1 _09203_ (.A(_01332_),
    .B(_01335_),
    .X(_01336_));
 sky130_fd_sc_hd__and2_1 _09204_ (.A(_01331_),
    .B(_01336_),
    .X(_01337_));
 sky130_fd_sc_hd__nor2_1 _09205_ (.A(_01331_),
    .B(_01336_),
    .Y(_01338_));
 sky130_fd_sc_hd__or2_1 _09206_ (.A(_01337_),
    .B(_01338_),
    .X(_01340_));
 sky130_fd_sc_hd__and3_1 _09207_ (.A(_01144_),
    .B(_01330_),
    .C(_01340_),
    .X(_01341_));
 sky130_fd_sc_hd__a21oi_1 _09208_ (.A1(_01144_),
    .A2(_01330_),
    .B1(_01340_),
    .Y(_01342_));
 sky130_fd_sc_hd__nor2_1 _09209_ (.A(_01341_),
    .B(_01342_),
    .Y(_01343_));
 sky130_fd_sc_hd__xnor2_1 _09210_ (.A(_01329_),
    .B(_01343_),
    .Y(_01344_));
 sky130_fd_sc_hd__nor2_1 _09211_ (.A(_01149_),
    .B(_01344_),
    .Y(_01345_));
 sky130_fd_sc_hd__and2_1 _09212_ (.A(_01149_),
    .B(_01344_),
    .X(_01346_));
 sky130_fd_sc_hd__nor2_1 _09213_ (.A(_01345_),
    .B(_01346_),
    .Y(_01347_));
 sky130_fd_sc_hd__xnor2_2 _09214_ (.A(_01316_),
    .B(_01347_),
    .Y(_01348_));
 sky130_fd_sc_hd__a21oi_1 _09215_ (.A1(_01155_),
    .A2(_01156_),
    .B1(_01154_),
    .Y(_01349_));
 sky130_fd_sc_hd__or2_2 _09216_ (.A(_01152_),
    .B(_01349_),
    .X(_01351_));
 sky130_fd_sc_hd__xor2_2 _09217_ (.A(_01348_),
    .B(_01351_),
    .X(_01352_));
 sky130_fd_sc_hd__xor2_1 _09218_ (.A(_01311_),
    .B(_01352_),
    .X(_01353_));
 sky130_fd_sc_hd__or2b_1 _09219_ (.A(_01310_),
    .B_N(_01352_),
    .X(_01354_));
 sky130_fd_sc_hd__a21bo_1 _09220_ (.A1(_01310_),
    .A2(_01353_),
    .B1_N(_01354_),
    .X(_01355_));
 sky130_fd_sc_hd__and3_2 _09221_ (.A(_01168_),
    .B(_01169_),
    .C(_01166_),
    .X(_01356_));
 sky130_fd_sc_hd__a21boi_1 _09222_ (.A1(_01168_),
    .A2(_01165_),
    .B1_N(_01162_),
    .Y(_01357_));
 sky130_fd_sc_hd__a21o_1 _09223_ (.A1(_00991_),
    .A2(_01356_),
    .B1(_01357_),
    .X(_01358_));
 sky130_fd_sc_hd__xnor2_2 _09224_ (.A(_01355_),
    .B(_01358_),
    .Y(_01359_));
 sky130_fd_sc_hd__o21a_1 _09225_ (.A1(_01057_),
    .A2(_01107_),
    .B1(_01110_),
    .X(_01360_));
 sky130_fd_sc_hd__a22oi_1 _09226_ (.A1(_00410_),
    .A2(_00376_),
    .B1(_00380_),
    .B2(_03015_),
    .Y(_01362_));
 sky130_fd_sc_hd__and3_1 _09227_ (.A(_00355_),
    .B(_02960_),
    .C(_04015_),
    .X(_01363_));
 sky130_fd_sc_hd__and2_1 _09228_ (.A(_04048_),
    .B(_01363_),
    .X(_01364_));
 sky130_fd_sc_hd__or2_1 _09229_ (.A(_01362_),
    .B(_01364_),
    .X(_01365_));
 sky130_fd_sc_hd__and2b_1 _09230_ (.A_N(_01071_),
    .B(_01079_),
    .X(_01366_));
 sky130_fd_sc_hd__a31oi_2 _09231_ (.A1(_01339_),
    .A2(_00604_),
    .A3(_01074_),
    .B1(_01073_),
    .Y(_01367_));
 sky130_fd_sc_hd__buf_2 _09232_ (.A(net47),
    .X(_01368_));
 sky130_fd_sc_hd__clkbuf_4 _09233_ (.A(_00959_),
    .X(_01369_));
 sky130_fd_sc_hd__a22oi_1 _09234_ (.A1(_04268_),
    .A2(_01368_),
    .B1(_01369_),
    .B2(_01372_),
    .Y(_01370_));
 sky130_fd_sc_hd__and4_1 _09235_ (.A(_01284_),
    .B(_01230_),
    .C(_01368_),
    .D(_00959_),
    .X(_01371_));
 sky130_fd_sc_hd__or2_1 _09236_ (.A(_01370_),
    .B(_01371_),
    .X(_01373_));
 sky130_fd_sc_hd__xor2_1 _09237_ (.A(_01367_),
    .B(_01373_),
    .X(_01374_));
 sky130_fd_sc_hd__and3_1 _09238_ (.A(_01072_),
    .B(_01078_),
    .C(_01374_),
    .X(_01375_));
 sky130_fd_sc_hd__a21oi_1 _09239_ (.A1(_01072_),
    .A2(_01078_),
    .B1(_01374_),
    .Y(_01376_));
 sky130_fd_sc_hd__nor2_1 _09240_ (.A(_01375_),
    .B(_01376_),
    .Y(_01377_));
 sky130_fd_sc_hd__o21a_1 _09241_ (.A1(_01366_),
    .A2(_01081_),
    .B1(_01377_),
    .X(_01378_));
 sky130_fd_sc_hd__nor3_1 _09242_ (.A(_01366_),
    .B(_01081_),
    .C(_01377_),
    .Y(_01379_));
 sky130_fd_sc_hd__nor2_1 _09243_ (.A(_01378_),
    .B(_01379_),
    .Y(_01380_));
 sky130_fd_sc_hd__and2b_1 _09244_ (.A_N(_01085_),
    .B(_01093_),
    .X(_01381_));
 sky130_fd_sc_hd__a31oi_2 _09245_ (.A1(_05566_),
    .A2(_00373_),
    .A3(_01089_),
    .B1(_01088_),
    .Y(_01382_));
 sky130_fd_sc_hd__a22oi_1 _09246_ (.A1(_03268_),
    .A2(_00612_),
    .B1(_00613_),
    .B2(_05577_),
    .Y(_01384_));
 sky130_fd_sc_hd__and4_2 _09247_ (.A(_02664_),
    .B(_02719_),
    .C(_00780_),
    .D(_00777_),
    .X(_01385_));
 sky130_fd_sc_hd__or2_1 _09248_ (.A(_01384_),
    .B(_01385_),
    .X(_01386_));
 sky130_fd_sc_hd__xor2_1 _09249_ (.A(_01382_),
    .B(_01386_),
    .X(_01387_));
 sky130_fd_sc_hd__and3_1 _09250_ (.A(_01086_),
    .B(_01092_),
    .C(_01387_),
    .X(_01388_));
 sky130_fd_sc_hd__a21oi_1 _09251_ (.A1(_01086_),
    .A2(_01092_),
    .B1(_01387_),
    .Y(_01389_));
 sky130_fd_sc_hd__nor2_1 _09252_ (.A(_01388_),
    .B(_01389_),
    .Y(_01390_));
 sky130_fd_sc_hd__o21a_1 _09253_ (.A1(_01381_),
    .A2(_01095_),
    .B1(_01390_),
    .X(_01391_));
 sky130_fd_sc_hd__nor3_1 _09254_ (.A(_01381_),
    .B(_01095_),
    .C(_01390_),
    .Y(_01392_));
 sky130_fd_sc_hd__nor2_1 _09255_ (.A(_01391_),
    .B(_01392_),
    .Y(_01393_));
 sky130_fd_sc_hd__xnor2_1 _09256_ (.A(_01380_),
    .B(_01393_),
    .Y(_01395_));
 sky130_fd_sc_hd__and2_1 _09257_ (.A(_01099_),
    .B(_01395_),
    .X(_01396_));
 sky130_fd_sc_hd__nor2_1 _09258_ (.A(_01099_),
    .B(_01395_),
    .Y(_01397_));
 sky130_fd_sc_hd__or2_1 _09259_ (.A(_01396_),
    .B(_01397_),
    .X(_01398_));
 sky130_fd_sc_hd__and3_1 _09260_ (.A(_02116_),
    .B(_02160_),
    .C(_00605_),
    .X(_01399_));
 sky130_fd_sc_hd__clkbuf_4 _09261_ (.A(_00608_),
    .X(_01400_));
 sky130_fd_sc_hd__a22o_1 _09262_ (.A1(_02171_),
    .A2(_00460_),
    .B1(_01400_),
    .B2(_02467_),
    .X(_01401_));
 sky130_fd_sc_hd__a21bo_1 _09263_ (.A1(_01066_),
    .A2(_01399_),
    .B1_N(_01401_),
    .X(_01402_));
 sky130_fd_sc_hd__xnor2_1 _09264_ (.A(_01398_),
    .B(_01402_),
    .Y(_01403_));
 sky130_fd_sc_hd__a21o_1 _09265_ (.A1(_01067_),
    .A2(_01103_),
    .B1(_01102_),
    .X(_01404_));
 sky130_fd_sc_hd__xor2_1 _09266_ (.A(_01403_),
    .B(_01404_),
    .X(_01406_));
 sky130_fd_sc_hd__and3_1 _09267_ (.A(_01064_),
    .B(_01105_),
    .C(_01406_),
    .X(_01407_));
 sky130_fd_sc_hd__a21oi_1 _09268_ (.A1(_01064_),
    .A2(_01105_),
    .B1(_01406_),
    .Y(_01408_));
 sky130_fd_sc_hd__or2_1 _09269_ (.A(_01407_),
    .B(_01408_),
    .X(_01409_));
 sky130_fd_sc_hd__clkbuf_4 _09270_ (.A(net50),
    .X(_01410_));
 sky130_fd_sc_hd__clkbuf_4 _09271_ (.A(_01410_),
    .X(_01411_));
 sky130_fd_sc_hd__clkbuf_4 _09272_ (.A(_01411_),
    .X(_01412_));
 sky130_fd_sc_hd__clkbuf_4 _09273_ (.A(_01412_),
    .X(_01413_));
 sky130_fd_sc_hd__clkbuf_4 _09274_ (.A(_01413_),
    .X(_01414_));
 sky130_fd_sc_hd__buf_4 _09275_ (.A(_01414_),
    .X(_01415_));
 sky130_fd_sc_hd__a22oi_1 _09276_ (.A1(_02051_),
    .A2(_01062_),
    .B1(_01415_),
    .B2(_00464_),
    .Y(_01417_));
 sky130_fd_sc_hd__and3_1 _09277_ (.A(_00431_),
    .B(_04169_),
    .C(net50),
    .X(_01418_));
 sky130_fd_sc_hd__and2_1 _09278_ (.A(_01058_),
    .B(_01418_),
    .X(_01419_));
 sky130_fd_sc_hd__or2_1 _09279_ (.A(_01417_),
    .B(_01419_),
    .X(_01420_));
 sky130_fd_sc_hd__xnor2_1 _09280_ (.A(_01409_),
    .B(_01420_),
    .Y(_01421_));
 sky130_fd_sc_hd__xor2_1 _09281_ (.A(_01365_),
    .B(_01421_),
    .X(_01422_));
 sky130_fd_sc_hd__and2_1 _09282_ (.A(_01360_),
    .B(_01422_),
    .X(_01423_));
 sky130_fd_sc_hd__nor2_1 _09283_ (.A(_01360_),
    .B(_01422_),
    .Y(_01424_));
 sky130_fd_sc_hd__nor2_1 _09284_ (.A(_01423_),
    .B(_01424_),
    .Y(_01425_));
 sky130_fd_sc_hd__xnor2_2 _09285_ (.A(_01359_),
    .B(_01425_),
    .Y(_01426_));
 sky130_fd_sc_hd__xnor2_4 _09286_ (.A(_01309_),
    .B(_01426_),
    .Y(_01428_));
 sky130_fd_sc_hd__nand2_1 _09287_ (.A(_01112_),
    .B(_01174_),
    .Y(_01429_));
 sky130_fd_sc_hd__nor2_1 _09288_ (.A(_01112_),
    .B(_01174_),
    .Y(_01430_));
 sky130_fd_sc_hd__a21oi_4 _09289_ (.A1(_01429_),
    .A2(_01233_),
    .B1(_01430_),
    .Y(_01431_));
 sky130_fd_sc_hd__xnor2_4 _09290_ (.A(_01428_),
    .B(_01431_),
    .Y(_01432_));
 sky130_fd_sc_hd__xnor2_4 _09291_ (.A(_01243_),
    .B(_01432_),
    .Y(_01433_));
 sky130_fd_sc_hd__or2_4 _09292_ (.A(_01054_),
    .B(_01239_),
    .X(_01434_));
 sky130_fd_sc_hd__nor2_1 _09293_ (.A(_00899_),
    .B(_01053_),
    .Y(_01435_));
 sky130_fd_sc_hd__o21a_1 _09294_ (.A1(_01056_),
    .A2(_01435_),
    .B1(_01238_),
    .X(_01436_));
 sky130_fd_sc_hd__o21bai_4 _09295_ (.A1(_00898_),
    .A2(_01434_),
    .B1_N(_01436_),
    .Y(_01437_));
 sky130_fd_sc_hd__xor2_4 _09296_ (.A(_01433_),
    .B(_01437_),
    .X(net82));
 sky130_fd_sc_hd__inv_2 _09297_ (.A(_01431_),
    .Y(_01439_));
 sky130_fd_sc_hd__or3b_2 _09298_ (.A(_01355_),
    .B(_01163_),
    .C_N(_01162_),
    .X(_01440_));
 sky130_fd_sc_hd__inv_2 _09299_ (.A(_01440_),
    .Y(_01441_));
 sky130_fd_sc_hd__a21oi_2 _09300_ (.A1(_01170_),
    .A2(_01171_),
    .B1(_01440_),
    .Y(_01442_));
 sky130_fd_sc_hd__a31oi_4 _09301_ (.A1(_00557_),
    .A2(_01167_),
    .A3(_01441_),
    .B1(_01442_),
    .Y(_01443_));
 sky130_fd_sc_hd__o21a_1 _09302_ (.A1(_01165_),
    .A2(_01353_),
    .B1(_01354_),
    .X(_01444_));
 sky130_fd_sc_hd__nor2_1 _09303_ (.A(_01348_),
    .B(_01351_),
    .Y(_01445_));
 sky130_fd_sc_hd__and2b_1 _09304_ (.A_N(_01311_),
    .B(_01352_),
    .X(_01446_));
 sky130_fd_sc_hd__nand2_1 _09305_ (.A(_01329_),
    .B(_01343_),
    .Y(_01447_));
 sky130_fd_sc_hd__and2b_1 _09306_ (.A_N(_01318_),
    .B(_01323_),
    .X(_01449_));
 sky130_fd_sc_hd__nor2_1 _09307_ (.A(_01319_),
    .B(_01322_),
    .Y(_01450_));
 sky130_fd_sc_hd__nand2_1 _09308_ (.A(_00844_),
    .B(_00819_),
    .Y(_01451_));
 sky130_fd_sc_hd__and3_1 _09309_ (.A(_00843_),
    .B(_00818_),
    .C(_01451_),
    .X(_01452_));
 sky130_fd_sc_hd__xor2_1 _09310_ (.A(_01450_),
    .B(_01452_),
    .X(_01453_));
 sky130_fd_sc_hd__nor3_1 _09311_ (.A(_01449_),
    .B(_01327_),
    .C(_01453_),
    .Y(_01454_));
 sky130_fd_sc_hd__o21a_1 _09312_ (.A1(_01449_),
    .A2(_01327_),
    .B1(_01453_),
    .X(_01455_));
 sky130_fd_sc_hd__nor2_1 _09313_ (.A(_01454_),
    .B(_01455_),
    .Y(_01456_));
 sky130_fd_sc_hd__nor2_1 _09314_ (.A(_01332_),
    .B(_01335_),
    .Y(_01457_));
 sky130_fd_sc_hd__and3_1 _09315_ (.A(_00262_),
    .B(_00859_),
    .C(_01136_),
    .X(_01458_));
 sky130_fd_sc_hd__xor2_1 _09316_ (.A(_01457_),
    .B(_01458_),
    .X(_01460_));
 sky130_fd_sc_hd__nor3_1 _09317_ (.A(_01337_),
    .B(_01342_),
    .C(_01460_),
    .Y(_01461_));
 sky130_fd_sc_hd__o21a_1 _09318_ (.A1(_01337_),
    .A2(_01342_),
    .B1(_01460_),
    .X(_01462_));
 sky130_fd_sc_hd__nor2_2 _09319_ (.A(_01461_),
    .B(_01462_),
    .Y(_01463_));
 sky130_fd_sc_hd__xnor2_1 _09320_ (.A(_01456_),
    .B(_01463_),
    .Y(_01464_));
 sky130_fd_sc_hd__nand2_1 _09321_ (.A(_01447_),
    .B(_01464_),
    .Y(_01465_));
 sky130_fd_sc_hd__or2_1 _09322_ (.A(_01447_),
    .B(_01464_),
    .X(_01466_));
 sky130_fd_sc_hd__and2_1 _09323_ (.A(_01465_),
    .B(_01466_),
    .X(_01467_));
 sky130_fd_sc_hd__and3_1 _09324_ (.A(_00844_),
    .B(_00654_),
    .C(_00635_),
    .X(_01468_));
 sky130_fd_sc_hd__a22o_1 _09325_ (.A1(_00654_),
    .A2(_00635_),
    .B1(_07040_),
    .B2(_00844_),
    .X(_01469_));
 sky130_fd_sc_hd__a21bo_1 _09326_ (.A1(_00526_),
    .A2(_01468_),
    .B1_N(_01469_),
    .X(_01471_));
 sky130_fd_sc_hd__clkbuf_4 _09327_ (.A(_00145_),
    .X(_01472_));
 sky130_fd_sc_hd__clkbuf_4 _09328_ (.A(_01472_),
    .X(_01473_));
 sky130_fd_sc_hd__nand2_1 _09329_ (.A(_00544_),
    .B(_01473_),
    .Y(_01474_));
 sky130_fd_sc_hd__xnor2_1 _09330_ (.A(_01471_),
    .B(_01474_),
    .Y(_01475_));
 sky130_fd_sc_hd__nor2_1 _09331_ (.A(_01315_),
    .B(_01475_),
    .Y(_01476_));
 sky130_fd_sc_hd__and2_1 _09332_ (.A(_01315_),
    .B(_01475_),
    .X(_01477_));
 sky130_fd_sc_hd__or2_1 _09333_ (.A(_01476_),
    .B(_01477_),
    .X(_01478_));
 sky130_fd_sc_hd__xnor2_1 _09334_ (.A(_01467_),
    .B(_01478_),
    .Y(_01479_));
 sky130_fd_sc_hd__inv_2 _09335_ (.A(_01346_),
    .Y(_01480_));
 sky130_fd_sc_hd__a21oi_1 _09336_ (.A1(_01316_),
    .A2(_01480_),
    .B1(_01345_),
    .Y(_01482_));
 sky130_fd_sc_hd__xnor2_1 _09337_ (.A(_01479_),
    .B(_01482_),
    .Y(_01483_));
 sky130_fd_sc_hd__or3_1 _09338_ (.A(_01445_),
    .B(_01446_),
    .C(_01483_),
    .X(_01484_));
 sky130_fd_sc_hd__o21ai_2 _09339_ (.A1(_01445_),
    .A2(_01446_),
    .B1(_01483_),
    .Y(_01485_));
 sky130_fd_sc_hd__nand2_2 _09340_ (.A(_01484_),
    .B(_01485_),
    .Y(_01486_));
 sky130_fd_sc_hd__a21o_1 _09341_ (.A1(_01443_),
    .A2(_01444_),
    .B1(_01486_),
    .X(_01487_));
 sky130_fd_sc_hd__inv_2 _09342_ (.A(_01444_),
    .Y(_01488_));
 sky130_fd_sc_hd__a31o_1 _09343_ (.A1(_00557_),
    .A2(_01167_),
    .A3(_01441_),
    .B1(_01442_),
    .X(_01489_));
 sky130_fd_sc_hd__or3b_1 _09344_ (.A(_01488_),
    .B(_01489_),
    .C_N(_01486_),
    .X(_01490_));
 sky130_fd_sc_hd__a21o_1 _09345_ (.A1(_01409_),
    .A2(_01420_),
    .B1(_01365_),
    .X(_01491_));
 sky130_fd_sc_hd__o21ai_1 _09346_ (.A1(_01409_),
    .A2(_01420_),
    .B1(_01491_),
    .Y(_01493_));
 sky130_fd_sc_hd__a22o_1 _09347_ (.A1(_02960_),
    .A2(_04015_),
    .B1(_04180_),
    .B2(_00355_),
    .X(_01494_));
 sky130_fd_sc_hd__a21bo_1 _09348_ (.A1(_00612_),
    .A2(_01363_),
    .B1_N(_01494_),
    .X(_01495_));
 sky130_fd_sc_hd__nand2_1 _09349_ (.A(_05192_),
    .B(net40),
    .Y(_01496_));
 sky130_fd_sc_hd__xor2_1 _09350_ (.A(_01495_),
    .B(_01496_),
    .X(_01497_));
 sky130_fd_sc_hd__and2_1 _09351_ (.A(_01364_),
    .B(_01497_),
    .X(_01498_));
 sky130_fd_sc_hd__nor2_1 _09352_ (.A(_01364_),
    .B(_01497_),
    .Y(_01499_));
 sky130_fd_sc_hd__or2_2 _09353_ (.A(_01498_),
    .B(_01499_),
    .X(_01500_));
 sky130_fd_sc_hd__nand2_1 _09354_ (.A(_01380_),
    .B(_01393_),
    .Y(_01501_));
 sky130_fd_sc_hd__nor2_1 _09355_ (.A(_01367_),
    .B(_01373_),
    .Y(_01502_));
 sky130_fd_sc_hd__clkbuf_4 _09356_ (.A(_01369_),
    .X(_01504_));
 sky130_fd_sc_hd__clkbuf_4 _09357_ (.A(_01504_),
    .X(_01505_));
 sky130_fd_sc_hd__buf_2 _09358_ (.A(_01368_),
    .X(_01506_));
 sky130_fd_sc_hd__clkbuf_4 _09359_ (.A(_01506_),
    .X(_01507_));
 sky130_fd_sc_hd__clkbuf_4 _09360_ (.A(_01507_),
    .X(_01508_));
 sky130_fd_sc_hd__nand2_1 _09361_ (.A(_01383_),
    .B(_01508_),
    .Y(_01509_));
 sky130_fd_sc_hd__and3_1 _09362_ (.A(_01350_),
    .B(_01505_),
    .C(_01509_),
    .X(_01510_));
 sky130_fd_sc_hd__xor2_1 _09363_ (.A(_01502_),
    .B(_01510_),
    .X(_01511_));
 sky130_fd_sc_hd__o21a_1 _09364_ (.A1(_01375_),
    .A2(_01378_),
    .B1(_01511_),
    .X(_01512_));
 sky130_fd_sc_hd__nor3_1 _09365_ (.A(_01375_),
    .B(_01378_),
    .C(_01511_),
    .Y(_01513_));
 sky130_fd_sc_hd__nor2_1 _09366_ (.A(_01512_),
    .B(_01513_),
    .Y(_01515_));
 sky130_fd_sc_hd__nor2_1 _09367_ (.A(_01382_),
    .B(_01386_),
    .Y(_01516_));
 sky130_fd_sc_hd__clkbuf_4 _09368_ (.A(_00779_),
    .X(_01517_));
 sky130_fd_sc_hd__clkbuf_4 _09369_ (.A(_00784_),
    .X(_01518_));
 sky130_fd_sc_hd__nand2_1 _09370_ (.A(_06461_),
    .B(_01518_),
    .Y(_01519_));
 sky130_fd_sc_hd__and3_2 _09371_ (.A(_06483_),
    .B(_01517_),
    .C(_01519_),
    .X(_01520_));
 sky130_fd_sc_hd__xor2_1 _09372_ (.A(_01516_),
    .B(_01520_),
    .X(_01521_));
 sky130_fd_sc_hd__o21a_1 _09373_ (.A1(_01388_),
    .A2(_01391_),
    .B1(_01521_),
    .X(_01522_));
 sky130_fd_sc_hd__nor3_1 _09374_ (.A(_01388_),
    .B(_01391_),
    .C(_01521_),
    .Y(_01523_));
 sky130_fd_sc_hd__nor2_1 _09375_ (.A(_01522_),
    .B(_01523_),
    .Y(_01524_));
 sky130_fd_sc_hd__xnor2_1 _09376_ (.A(_01515_),
    .B(_01524_),
    .Y(_01526_));
 sky130_fd_sc_hd__nor2_1 _09377_ (.A(_01501_),
    .B(_01526_),
    .Y(_01527_));
 sky130_fd_sc_hd__and2_1 _09378_ (.A(_01501_),
    .B(_01526_),
    .X(_01528_));
 sky130_fd_sc_hd__nor2_1 _09379_ (.A(_01527_),
    .B(_01528_),
    .Y(_01529_));
 sky130_fd_sc_hd__a22o_1 _09380_ (.A1(_02160_),
    .A2(_00605_),
    .B1(_01508_),
    .B2(_02116_),
    .X(_01530_));
 sky130_fd_sc_hd__nand2_1 _09381_ (.A(_01508_),
    .B(_01399_),
    .Y(_01531_));
 sky130_fd_sc_hd__nand2_1 _09382_ (.A(_01530_),
    .B(_01531_),
    .Y(_01532_));
 sky130_fd_sc_hd__nand2_1 _09383_ (.A(_06472_),
    .B(_00458_),
    .Y(_01533_));
 sky130_fd_sc_hd__xor2_1 _09384_ (.A(_01532_),
    .B(_01533_),
    .X(_01534_));
 sky130_fd_sc_hd__and3_1 _09385_ (.A(_00459_),
    .B(_01399_),
    .C(_01534_),
    .X(_01535_));
 sky130_fd_sc_hd__a21oi_1 _09386_ (.A1(_00460_),
    .A2(_01399_),
    .B1(_01534_),
    .Y(_01537_));
 sky130_fd_sc_hd__or2_1 _09387_ (.A(_01535_),
    .B(_01537_),
    .X(_01538_));
 sky130_fd_sc_hd__xnor2_2 _09388_ (.A(_01529_),
    .B(_01538_),
    .Y(_01539_));
 sky130_fd_sc_hd__o21ba_1 _09389_ (.A1(_01396_),
    .A2(_01402_),
    .B1_N(_01397_),
    .X(_01540_));
 sky130_fd_sc_hd__xnor2_2 _09390_ (.A(_01539_),
    .B(_01540_),
    .Y(_01541_));
 sky130_fd_sc_hd__nor2_1 _09391_ (.A(_01403_),
    .B(_01404_),
    .Y(_01542_));
 sky130_fd_sc_hd__a31o_1 _09392_ (.A1(_01064_),
    .A2(_01105_),
    .A3(_01406_),
    .B1(_01542_),
    .X(_01543_));
 sky130_fd_sc_hd__xnor2_2 _09393_ (.A(_01541_),
    .B(_01543_),
    .Y(_01544_));
 sky130_fd_sc_hd__buf_2 _09394_ (.A(net51),
    .X(_01545_));
 sky130_fd_sc_hd__buf_2 _09395_ (.A(_01545_),
    .X(_01546_));
 sky130_fd_sc_hd__a22o_1 _09396_ (.A1(_04169_),
    .A2(net50),
    .B1(_01545_),
    .B2(_00431_),
    .X(_01548_));
 sky130_fd_sc_hd__a21bo_1 _09397_ (.A1(_01546_),
    .A2(_01418_),
    .B1_N(_01548_),
    .X(_01549_));
 sky130_fd_sc_hd__nand2_1 _09398_ (.A(_01372_),
    .B(net49),
    .Y(_01550_));
 sky130_fd_sc_hd__xor2_1 _09399_ (.A(_01549_),
    .B(_01550_),
    .X(_01551_));
 sky130_fd_sc_hd__and2_1 _09400_ (.A(_01419_),
    .B(_01551_),
    .X(_01552_));
 sky130_fd_sc_hd__nor2_1 _09401_ (.A(_01419_),
    .B(_01551_),
    .Y(_01553_));
 sky130_fd_sc_hd__or2_1 _09402_ (.A(_01552_),
    .B(_01553_),
    .X(_01554_));
 sky130_fd_sc_hd__xor2_1 _09403_ (.A(_01544_),
    .B(_01554_),
    .X(_01555_));
 sky130_fd_sc_hd__xnor2_1 _09404_ (.A(_01500_),
    .B(_01555_),
    .Y(_01556_));
 sky130_fd_sc_hd__xor2_1 _09405_ (.A(_01493_),
    .B(_01556_),
    .X(_01557_));
 sky130_fd_sc_hd__xor2_1 _09406_ (.A(_01423_),
    .B(_01557_),
    .X(_01559_));
 sky130_fd_sc_hd__a21oi_1 _09407_ (.A1(_01487_),
    .A2(_01490_),
    .B1(_01559_),
    .Y(_01560_));
 sky130_fd_sc_hd__and3_1 _09408_ (.A(_01559_),
    .B(_01487_),
    .C(_01490_),
    .X(_01561_));
 sky130_fd_sc_hd__o21ai_1 _09409_ (.A1(_01298_),
    .A2(_01299_),
    .B1(_01303_),
    .Y(_01562_));
 sky130_fd_sc_hd__a32o_2 _09410_ (.A1(_01300_),
    .A2(_01301_),
    .A3(_01302_),
    .B1(_01562_),
    .B2(_01256_),
    .X(_01563_));
 sky130_fd_sc_hd__buf_2 _09411_ (.A(net19),
    .X(_01564_));
 sky130_fd_sc_hd__a22o_1 _09412_ (.A1(_04510_),
    .A2(_01177_),
    .B1(_01246_),
    .B2(_00661_),
    .X(_01565_));
 sky130_fd_sc_hd__inv_2 _09413_ (.A(_01565_),
    .Y(_01566_));
 sky130_fd_sc_hd__and4_1 _09414_ (.A(_04510_),
    .B(_00661_),
    .C(net17),
    .D(net18),
    .X(_01567_));
 sky130_fd_sc_hd__o2bb2a_1 _09415_ (.A1_N(_00322_),
    .A2_N(_01564_),
    .B1(_01566_),
    .B2(_01567_),
    .X(_01568_));
 sky130_fd_sc_hd__and4b_1 _09416_ (.A_N(_01567_),
    .B(_01564_),
    .C(_00311_),
    .D(_01565_),
    .X(_01570_));
 sky130_fd_sc_hd__or2_2 _09417_ (.A(_01568_),
    .B(_01570_),
    .X(_01571_));
 sky130_fd_sc_hd__xnor2_4 _09418_ (.A(_01255_),
    .B(_01571_),
    .Y(_01572_));
 sky130_fd_sc_hd__nand2_1 _09419_ (.A(_01269_),
    .B(_01282_),
    .Y(_01573_));
 sky130_fd_sc_hd__and3_1 _09420_ (.A(_01193_),
    .B(_01199_),
    .C(_01265_),
    .X(_01574_));
 sky130_fd_sc_hd__nand2_1 _09421_ (.A(_00138_),
    .B(_00742_),
    .Y(_01575_));
 sky130_fd_sc_hd__nand4_1 _09422_ (.A(_06428_),
    .B(_00745_),
    .C(_01575_),
    .D(_01263_),
    .Y(_01576_));
 sky130_fd_sc_hd__a31o_1 _09423_ (.A1(_06417_),
    .A2(_00745_),
    .A3(_01575_),
    .B1(_01263_),
    .X(_01577_));
 sky130_fd_sc_hd__and2_1 _09424_ (.A(_01576_),
    .B(_01577_),
    .X(_01578_));
 sky130_fd_sc_hd__o21ai_1 _09425_ (.A1(_01574_),
    .A2(_01267_),
    .B1(_01578_),
    .Y(_01579_));
 sky130_fd_sc_hd__or3_1 _09426_ (.A(_01574_),
    .B(_01267_),
    .C(_01578_),
    .X(_01581_));
 sky130_fd_sc_hd__and2_1 _09427_ (.A(_01579_),
    .B(_01581_),
    .X(_01582_));
 sky130_fd_sc_hd__and3_1 _09428_ (.A(_01207_),
    .B(_01214_),
    .C(_01278_),
    .X(_01583_));
 sky130_fd_sc_hd__buf_4 _09429_ (.A(_01211_),
    .X(_01584_));
 sky130_fd_sc_hd__buf_4 _09430_ (.A(_01584_),
    .X(_01585_));
 sky130_fd_sc_hd__buf_4 _09431_ (.A(_01272_),
    .X(_01586_));
 sky130_fd_sc_hd__nand2_1 _09432_ (.A(_00159_),
    .B(_01586_),
    .Y(_01587_));
 sky130_fd_sc_hd__nand4_1 _09433_ (.A(_00157_),
    .B(_01585_),
    .C(_01587_),
    .D(_01276_),
    .Y(_01588_));
 sky130_fd_sc_hd__a31o_1 _09434_ (.A1(_00157_),
    .A2(_01584_),
    .A3(_01587_),
    .B1(_01276_),
    .X(_01589_));
 sky130_fd_sc_hd__and2_1 _09435_ (.A(_01588_),
    .B(_01589_),
    .X(_01590_));
 sky130_fd_sc_hd__o21ai_1 _09436_ (.A1(_01583_),
    .A2(_01280_),
    .B1(_01590_),
    .Y(_01592_));
 sky130_fd_sc_hd__or3_1 _09437_ (.A(_01583_),
    .B(_01280_),
    .C(_01590_),
    .X(_01593_));
 sky130_fd_sc_hd__and2_1 _09438_ (.A(_01592_),
    .B(_01593_),
    .X(_01594_));
 sky130_fd_sc_hd__xnor2_1 _09439_ (.A(_01582_),
    .B(_01594_),
    .Y(_01595_));
 sky130_fd_sc_hd__xnor2_1 _09440_ (.A(_01573_),
    .B(_01595_),
    .Y(_01596_));
 sky130_fd_sc_hd__and3_1 _09441_ (.A(_06439_),
    .B(_02018_),
    .C(_00574_),
    .X(_01597_));
 sky130_fd_sc_hd__a22o_1 _09442_ (.A1(_06439_),
    .A2(_00414_),
    .B1(_00574_),
    .B2(_02018_),
    .X(_01598_));
 sky130_fd_sc_hd__a21bo_1 _09443_ (.A1(_00416_),
    .A2(_01597_),
    .B1_N(_01598_),
    .X(_01599_));
 sky130_fd_sc_hd__clkbuf_4 _09444_ (.A(_01586_),
    .X(_01600_));
 sky130_fd_sc_hd__clkbuf_4 _09445_ (.A(_01600_),
    .X(_01601_));
 sky130_fd_sc_hd__nand2_1 _09446_ (.A(_02335_),
    .B(_01601_),
    .Y(_01603_));
 sky130_fd_sc_hd__xnor2_1 _09447_ (.A(_01599_),
    .B(_01603_),
    .Y(_01604_));
 sky130_fd_sc_hd__nor2_1 _09448_ (.A(_01292_),
    .B(_01604_),
    .Y(_01605_));
 sky130_fd_sc_hd__and2_1 _09449_ (.A(_01292_),
    .B(_01604_),
    .X(_01606_));
 sky130_fd_sc_hd__or2_2 _09450_ (.A(_01605_),
    .B(_01606_),
    .X(_01607_));
 sky130_fd_sc_hd__xnor2_2 _09451_ (.A(_01596_),
    .B(_01607_),
    .Y(_01608_));
 sky130_fd_sc_hd__a21bo_1 _09452_ (.A1(_01285_),
    .A2(_01293_),
    .B1_N(_01286_),
    .X(_01609_));
 sky130_fd_sc_hd__xnor2_2 _09453_ (.A(_01608_),
    .B(_01609_),
    .Y(_01610_));
 sky130_fd_sc_hd__and2b_1 _09454_ (.A_N(_01296_),
    .B(_01294_),
    .X(_01611_));
 sky130_fd_sc_hd__a31o_4 _09455_ (.A1(_01187_),
    .A2(_01227_),
    .A3(_01297_),
    .B1(_01611_),
    .X(_01612_));
 sky130_fd_sc_hd__xnor2_2 _09456_ (.A(_01610_),
    .B(_01612_),
    .Y(_01614_));
 sky130_fd_sc_hd__a22o_1 _09457_ (.A1(_06820_),
    .A2(net8),
    .B1(net9),
    .B2(net64),
    .X(_01615_));
 sky130_fd_sc_hd__inv_2 _09458_ (.A(_01615_),
    .Y(_01616_));
 sky130_fd_sc_hd__and4_1 _09459_ (.A(net64),
    .B(_06820_),
    .C(net8),
    .D(net9),
    .X(_01617_));
 sky130_fd_sc_hd__o2bb2a_1 _09460_ (.A1_N(_00475_),
    .A2_N(_03894_),
    .B1(_01616_),
    .B2(_01617_),
    .X(_01618_));
 sky130_fd_sc_hd__and4b_1 _09461_ (.A_N(_01617_),
    .B(_03894_),
    .C(_00475_),
    .D(_01615_),
    .X(_01619_));
 sky130_fd_sc_hd__or2_2 _09462_ (.A(_01618_),
    .B(_01619_),
    .X(_01620_));
 sky130_fd_sc_hd__xnor2_2 _09463_ (.A(_01302_),
    .B(_01620_),
    .Y(_01621_));
 sky130_fd_sc_hd__xor2_2 _09464_ (.A(_01614_),
    .B(_01621_),
    .X(_01622_));
 sky130_fd_sc_hd__xnor2_4 _09465_ (.A(_01572_),
    .B(_01622_),
    .Y(_01623_));
 sky130_fd_sc_hd__xor2_4 _09466_ (.A(_01563_),
    .B(_01623_),
    .X(_01625_));
 sky130_fd_sc_hd__xor2_4 _09467_ (.A(_01307_),
    .B(_01625_),
    .X(_01626_));
 sky130_fd_sc_hd__o21a_1 _09468_ (.A1(_01560_),
    .A2(_01561_),
    .B1(_01626_),
    .X(_01627_));
 sky130_fd_sc_hd__nor3_1 _09469_ (.A(_01626_),
    .B(_01560_),
    .C(_01561_),
    .Y(_01628_));
 sky130_fd_sc_hd__or2_1 _09470_ (.A(_01359_),
    .B(_01425_),
    .X(_01629_));
 sky130_fd_sc_hd__a21o_1 _09471_ (.A1(_01359_),
    .A2(_01425_),
    .B1(_01309_),
    .X(_01630_));
 sky130_fd_sc_hd__o211a_1 _09472_ (.A1(_01627_),
    .A2(_01628_),
    .B1(_01629_),
    .C1(_01630_),
    .X(_01631_));
 sky130_fd_sc_hd__a211oi_2 _09473_ (.A1(_01629_),
    .A2(_01630_),
    .B1(_01627_),
    .C1(_01628_),
    .Y(_01632_));
 sky130_fd_sc_hd__or4b_4 _09474_ (.A(_01439_),
    .B(_01631_),
    .C(_01632_),
    .D_N(_01428_),
    .X(_01633_));
 sky130_fd_sc_hd__a2bb2o_1 _09475_ (.A1_N(_01631_),
    .A2_N(_01632_),
    .B1(_01428_),
    .B2(_01431_),
    .X(_01634_));
 sky130_fd_sc_hd__and2_4 _09476_ (.A(_01633_),
    .B(_01634_),
    .X(_01636_));
 sky130_fd_sc_hd__inv_2 _09477_ (.A(_01239_),
    .Y(_01637_));
 sky130_fd_sc_hd__a21oi_1 _09478_ (.A1(_01056_),
    .A2(_01238_),
    .B1(_01243_),
    .Y(_01638_));
 sky130_fd_sc_hd__nor2_1 _09479_ (.A(_01432_),
    .B(_01638_),
    .Y(_01639_));
 sky130_fd_sc_hd__a31o_2 _09480_ (.A1(_01637_),
    .A2(net131),
    .A3(_01433_),
    .B1(_01639_),
    .X(_01640_));
 sky130_fd_sc_hd__xor2_4 _09481_ (.A(_01636_),
    .B(_01640_),
    .X(net83));
 sky130_fd_sc_hd__inv_2 _09482_ (.A(_01243_),
    .Y(_01641_));
 sky130_fd_sc_hd__nand2_1 _09483_ (.A(_01428_),
    .B(_01431_),
    .Y(_01642_));
 sky130_fd_sc_hd__o21ai_2 _09484_ (.A1(_01641_),
    .A2(_01432_),
    .B1(_01642_),
    .Y(_01643_));
 sky130_fd_sc_hd__or2_1 _09485_ (.A(_01631_),
    .B(_01632_),
    .X(_01644_));
 sky130_fd_sc_hd__inv_2 _09486_ (.A(_01644_),
    .Y(_01646_));
 sky130_fd_sc_hd__a32oi_4 _09487_ (.A1(_01433_),
    .A2(_01436_),
    .A3(_01636_),
    .B1(_01643_),
    .B2(_01646_),
    .Y(_01647_));
 sky130_fd_sc_hd__or4bb_4 _09488_ (.A(_01434_),
    .B(_00898_),
    .C_N(_01433_),
    .D_N(_01636_),
    .X(_01648_));
 sky130_fd_sc_hd__nand2_2 _09489_ (.A(_01647_),
    .B(_01648_),
    .Y(_01649_));
 sky130_fd_sc_hd__a22oi_1 _09490_ (.A1(_03587_),
    .A2(_01545_),
    .B1(net52),
    .B2(_03576_),
    .Y(_01650_));
 sky130_fd_sc_hd__and4_1 _09491_ (.A(_00431_),
    .B(_04169_),
    .C(net51),
    .D(net52),
    .X(_01651_));
 sky130_fd_sc_hd__nor2_1 _09492_ (.A(_01650_),
    .B(_01651_),
    .Y(_01652_));
 sky130_fd_sc_hd__nand2_1 _09493_ (.A(_01372_),
    .B(net50),
    .Y(_01653_));
 sky130_fd_sc_hd__xor2_1 _09494_ (.A(_01652_),
    .B(_01653_),
    .X(_01654_));
 sky130_fd_sc_hd__and4_1 _09495_ (.A(_00431_),
    .B(_04169_),
    .C(net50),
    .D(net51),
    .X(_01655_));
 sky130_fd_sc_hd__a31o_1 _09496_ (.A1(_01284_),
    .A2(net49),
    .A3(_01548_),
    .B1(_01655_),
    .X(_01657_));
 sky130_fd_sc_hd__nand2_1 _09497_ (.A(_04268_),
    .B(net49),
    .Y(_01658_));
 sky130_fd_sc_hd__xor2_1 _09498_ (.A(_01657_),
    .B(_01658_),
    .X(_01659_));
 sky130_fd_sc_hd__xor2_1 _09499_ (.A(_01654_),
    .B(_01659_),
    .X(_01660_));
 sky130_fd_sc_hd__and2_1 _09500_ (.A(_01552_),
    .B(_01660_),
    .X(_01661_));
 sky130_fd_sc_hd__nor2_1 _09501_ (.A(_01552_),
    .B(_01660_),
    .Y(_01662_));
 sky130_fd_sc_hd__or2_1 _09502_ (.A(_01661_),
    .B(_01662_),
    .X(_01663_));
 sky130_fd_sc_hd__clkbuf_4 _09503_ (.A(_01508_),
    .X(_01664_));
 sky130_fd_sc_hd__a22oi_2 _09504_ (.A1(_02160_),
    .A2(_01664_),
    .B1(_01505_),
    .B2(_02116_),
    .Y(_01665_));
 sky130_fd_sc_hd__and4_1 _09505_ (.A(_02116_),
    .B(_02160_),
    .C(_01508_),
    .D(_01504_),
    .X(_01666_));
 sky130_fd_sc_hd__or2_1 _09506_ (.A(_01665_),
    .B(_01666_),
    .X(_01668_));
 sky130_fd_sc_hd__nand2_1 _09507_ (.A(_06472_),
    .B(_00607_),
    .Y(_01669_));
 sky130_fd_sc_hd__xnor2_1 _09508_ (.A(_01668_),
    .B(_01669_),
    .Y(_01670_));
 sky130_fd_sc_hd__o21ai_1 _09509_ (.A1(_01532_),
    .A2(_01533_),
    .B1(_01531_),
    .Y(_01671_));
 sky130_fd_sc_hd__and3_1 _09510_ (.A(_06494_),
    .B(_00458_),
    .C(_01671_),
    .X(_01672_));
 sky130_fd_sc_hd__a21oi_1 _09511_ (.A1(_06494_),
    .A2(_00459_),
    .B1(_01671_),
    .Y(_01673_));
 sky130_fd_sc_hd__nor3_1 _09512_ (.A(_01670_),
    .B(_01672_),
    .C(_01673_),
    .Y(_01674_));
 sky130_fd_sc_hd__o21a_1 _09513_ (.A1(_01672_),
    .A2(_01673_),
    .B1(_01670_),
    .X(_01675_));
 sky130_fd_sc_hd__nor2_1 _09514_ (.A(_01674_),
    .B(_01675_),
    .Y(_01676_));
 sky130_fd_sc_hd__nand2_1 _09515_ (.A(_01535_),
    .B(_01676_),
    .Y(_01677_));
 sky130_fd_sc_hd__or2_1 _09516_ (.A(_01535_),
    .B(_01676_),
    .X(_01679_));
 sky130_fd_sc_hd__nand2_1 _09517_ (.A(_01677_),
    .B(_01679_),
    .Y(_01680_));
 sky130_fd_sc_hd__nand2_1 _09518_ (.A(_01515_),
    .B(_01524_),
    .Y(_01681_));
 sky130_fd_sc_hd__a211oi_2 _09519_ (.A1(_01502_),
    .A2(_01510_),
    .B1(_01512_),
    .C1(_01371_),
    .Y(_01682_));
 sky130_fd_sc_hd__a211oi_4 _09520_ (.A1(_01516_),
    .A2(_01520_),
    .B1(_01522_),
    .C1(_01385_),
    .Y(_01683_));
 sky130_fd_sc_hd__xnor2_2 _09521_ (.A(_01682_),
    .B(_01683_),
    .Y(_01684_));
 sky130_fd_sc_hd__xor2_1 _09522_ (.A(_01681_),
    .B(_01684_),
    .X(_01685_));
 sky130_fd_sc_hd__xnor2_1 _09523_ (.A(_01680_),
    .B(_01685_),
    .Y(_01686_));
 sky130_fd_sc_hd__o21a_1 _09524_ (.A1(_01501_),
    .A2(_01526_),
    .B1(_01538_),
    .X(_01687_));
 sky130_fd_sc_hd__or2_1 _09525_ (.A(_01528_),
    .B(_01687_),
    .X(_01688_));
 sky130_fd_sc_hd__and2b_1 _09526_ (.A_N(_01686_),
    .B(_01688_),
    .X(_01690_));
 sky130_fd_sc_hd__and2b_1 _09527_ (.A_N(_01688_),
    .B(_01686_),
    .X(_01691_));
 sky130_fd_sc_hd__nor2_1 _09528_ (.A(_01690_),
    .B(_01691_),
    .Y(_01692_));
 sky130_fd_sc_hd__inv_2 _09529_ (.A(_01540_),
    .Y(_01693_));
 sky130_fd_sc_hd__and2_1 _09530_ (.A(_01539_),
    .B(_01693_),
    .X(_01694_));
 sky130_fd_sc_hd__a21o_1 _09531_ (.A1(_01541_),
    .A2(_01543_),
    .B1(_01694_),
    .X(_01695_));
 sky130_fd_sc_hd__xnor2_2 _09532_ (.A(_01692_),
    .B(_01695_),
    .Y(_01696_));
 sky130_fd_sc_hd__xnor2_1 _09533_ (.A(_01663_),
    .B(_01696_),
    .Y(_01697_));
 sky130_fd_sc_hd__a22oi_1 _09534_ (.A1(_02971_),
    .A2(_04103_),
    .B1(_00777_),
    .B2(_00366_),
    .Y(_01698_));
 sky130_fd_sc_hd__and4_1 _09535_ (.A(_00355_),
    .B(_02960_),
    .C(_04180_),
    .D(_04191_),
    .X(_01699_));
 sky130_fd_sc_hd__nor2_1 _09536_ (.A(_01698_),
    .B(_01699_),
    .Y(_01701_));
 sky130_fd_sc_hd__nand2_1 _09537_ (.A(_05192_),
    .B(_04026_),
    .Y(_01702_));
 sky130_fd_sc_hd__xor2_1 _09538_ (.A(_01701_),
    .B(_01702_),
    .X(_01703_));
 sky130_fd_sc_hd__and4_1 _09539_ (.A(_00355_),
    .B(_02960_),
    .C(net41),
    .D(_04180_),
    .X(_01704_));
 sky130_fd_sc_hd__a31o_1 _09540_ (.A1(_05192_),
    .A2(net40),
    .A3(_01494_),
    .B1(_01704_),
    .X(_01705_));
 sky130_fd_sc_hd__nand2_1 _09541_ (.A(_04598_),
    .B(net40),
    .Y(_01706_));
 sky130_fd_sc_hd__xor2_1 _09542_ (.A(_01705_),
    .B(_01706_),
    .X(_01707_));
 sky130_fd_sc_hd__xor2_1 _09543_ (.A(_01703_),
    .B(_01707_),
    .X(_01708_));
 sky130_fd_sc_hd__and2_1 _09544_ (.A(_01498_),
    .B(_01708_),
    .X(_01709_));
 sky130_fd_sc_hd__nor2_1 _09545_ (.A(_01498_),
    .B(_01708_),
    .Y(_01710_));
 sky130_fd_sc_hd__or2_2 _09546_ (.A(_01709_),
    .B(_01710_),
    .X(_01712_));
 sky130_fd_sc_hd__xnor2_2 _09547_ (.A(_01697_),
    .B(_01712_),
    .Y(_01713_));
 sky130_fd_sc_hd__o21a_1 _09548_ (.A1(_01544_),
    .A2(_01554_),
    .B1(_01500_),
    .X(_01714_));
 sky130_fd_sc_hd__a21o_1 _09549_ (.A1(_01544_),
    .A2(_01554_),
    .B1(_01714_),
    .X(_01715_));
 sky130_fd_sc_hd__xor2_2 _09550_ (.A(_01713_),
    .B(_01715_),
    .X(_01716_));
 sky130_fd_sc_hd__a32o_1 _09551_ (.A1(_01360_),
    .A2(_01422_),
    .A3(_01557_),
    .B1(_01556_),
    .B2(_01493_),
    .X(_01717_));
 sky130_fd_sc_hd__xor2_1 _09552_ (.A(_01716_),
    .B(_01717_),
    .X(_01718_));
 sky130_fd_sc_hd__inv_2 _09553_ (.A(_01482_),
    .Y(_01719_));
 sky130_fd_sc_hd__nand2_1 _09554_ (.A(_01479_),
    .B(_01719_),
    .Y(_01720_));
 sky130_fd_sc_hd__nand2_1 _09555_ (.A(_01720_),
    .B(_01485_),
    .Y(_01721_));
 sky130_fd_sc_hd__nand2_1 _09556_ (.A(_01466_),
    .B(_01478_),
    .Y(_01723_));
 sky130_fd_sc_hd__and4_1 _09557_ (.A(_00843_),
    .B(_00844_),
    .C(_00635_),
    .D(_07040_),
    .X(_01724_));
 sky130_fd_sc_hd__a22oi_1 _09558_ (.A1(_00844_),
    .A2(_00635_),
    .B1(_07040_),
    .B2(_00843_),
    .Y(_01725_));
 sky130_fd_sc_hd__and4bb_1 _09559_ (.A_N(_01724_),
    .B_N(_01725_),
    .C(_00654_),
    .D(_01472_),
    .X(_01726_));
 sky130_fd_sc_hd__o2bb2a_1 _09560_ (.A1_N(_00654_),
    .A2_N(_01472_),
    .B1(_01724_),
    .B2(_01725_),
    .X(_01727_));
 sky130_fd_sc_hd__a32o_1 _09561_ (.A1(_00543_),
    .A2(_01472_),
    .A3(_01469_),
    .B1(_01468_),
    .B2(_07040_),
    .X(_01728_));
 sky130_fd_sc_hd__and3_1 _09562_ (.A(_00543_),
    .B(_00859_),
    .C(_01728_),
    .X(_01729_));
 sky130_fd_sc_hd__a21oi_1 _09563_ (.A1(_00544_),
    .A2(_00859_),
    .B1(_01728_),
    .Y(_01730_));
 sky130_fd_sc_hd__nor4_1 _09564_ (.A(_01726_),
    .B(_01727_),
    .C(_01729_),
    .D(_01730_),
    .Y(_01731_));
 sky130_fd_sc_hd__o22a_1 _09565_ (.A1(_01726_),
    .A2(_01727_),
    .B1(_01729_),
    .B2(_01730_),
    .X(_01732_));
 sky130_fd_sc_hd__nor2_1 _09566_ (.A(_01731_),
    .B(_01732_),
    .Y(_01734_));
 sky130_fd_sc_hd__nand2_1 _09567_ (.A(_01476_),
    .B(_01734_),
    .Y(_01735_));
 sky130_fd_sc_hd__or2_1 _09568_ (.A(_01476_),
    .B(_01734_),
    .X(_01736_));
 sky130_fd_sc_hd__and2_1 _09569_ (.A(_01735_),
    .B(_01736_),
    .X(_01737_));
 sky130_fd_sc_hd__nand2_1 _09570_ (.A(_01456_),
    .B(_01463_),
    .Y(_01738_));
 sky130_fd_sc_hd__a21o_1 _09571_ (.A1(_01450_),
    .A2(_01452_),
    .B1(_01455_),
    .X(_01739_));
 sky130_fd_sc_hd__and2b_1 _09572_ (.A_N(_01739_),
    .B(_01321_),
    .X(_01740_));
 sky130_fd_sc_hd__a211oi_4 _09573_ (.A1(_01457_),
    .A2(_01458_),
    .B1(_01462_),
    .C1(_01334_),
    .Y(_01741_));
 sky130_fd_sc_hd__xnor2_1 _09574_ (.A(_01740_),
    .B(_01741_),
    .Y(_01742_));
 sky130_fd_sc_hd__nand2_1 _09575_ (.A(_01738_),
    .B(_01742_),
    .Y(_01743_));
 sky130_fd_sc_hd__inv_2 _09576_ (.A(_01743_),
    .Y(_01745_));
 sky130_fd_sc_hd__nor2_1 _09577_ (.A(_01738_),
    .B(_01742_),
    .Y(_01746_));
 sky130_fd_sc_hd__nor2_1 _09578_ (.A(_01745_),
    .B(_01746_),
    .Y(_01747_));
 sky130_fd_sc_hd__xor2_1 _09579_ (.A(_01737_),
    .B(_01747_),
    .X(_01748_));
 sky130_fd_sc_hd__a21oi_1 _09580_ (.A1(_01465_),
    .A2(_01723_),
    .B1(_01748_),
    .Y(_01749_));
 sky130_fd_sc_hd__nand3_1 _09581_ (.A(_01465_),
    .B(_01723_),
    .C(_01748_),
    .Y(_01750_));
 sky130_fd_sc_hd__and2b_1 _09582_ (.A_N(_01749_),
    .B(_01750_),
    .X(_01751_));
 sky130_fd_sc_hd__xor2_2 _09583_ (.A(_01721_),
    .B(_01751_),
    .X(_01752_));
 sky130_fd_sc_hd__or2b_1 _09584_ (.A(_01486_),
    .B_N(_01752_),
    .X(_01753_));
 sky130_fd_sc_hd__a21o_1 _09585_ (.A1(_01443_),
    .A2(_01444_),
    .B1(_01753_),
    .X(_01754_));
 sky130_fd_sc_hd__nor2_2 _09586_ (.A(_01355_),
    .B(_01486_),
    .Y(_01756_));
 sky130_fd_sc_hd__a2bb2o_1 _09587_ (.A1_N(_01354_),
    .A2_N(_01486_),
    .B1(_01756_),
    .B2(_01357_),
    .X(_01757_));
 sky130_fd_sc_hd__a311o_1 _09588_ (.A1(_00991_),
    .A2(_01356_),
    .A3(_01756_),
    .B1(_01757_),
    .C1(_01752_),
    .X(_01758_));
 sky130_fd_sc_hd__and3_1 _09589_ (.A(_01718_),
    .B(_01754_),
    .C(_01758_),
    .X(_01759_));
 sky130_fd_sc_hd__a21oi_2 _09590_ (.A1(_01754_),
    .A2(_01758_),
    .B1(_01718_),
    .Y(_01760_));
 sky130_fd_sc_hd__and3_1 _09591_ (.A(_06818_),
    .B(_06820_),
    .C(net9),
    .X(_01761_));
 sky130_fd_sc_hd__a22o_1 _09592_ (.A1(_06818_),
    .A2(net8),
    .B1(net9),
    .B2(_06820_),
    .X(_01762_));
 sky130_fd_sc_hd__a21bo_1 _09593_ (.A1(_03685_),
    .A2(_01761_),
    .B1_N(_01762_),
    .X(_01763_));
 sky130_fd_sc_hd__nand2_1 _09594_ (.A(_03510_),
    .B(_03762_),
    .Y(_01764_));
 sky130_fd_sc_hd__xor2_1 _09595_ (.A(_01763_),
    .B(_01764_),
    .X(_01765_));
 sky130_fd_sc_hd__a31o_1 _09596_ (.A1(_00475_),
    .A2(net10),
    .A3(_01615_),
    .B1(_01617_),
    .X(_01767_));
 sky130_fd_sc_hd__nand2_1 _09597_ (.A(_00475_),
    .B(net11),
    .Y(_01768_));
 sky130_fd_sc_hd__xnor2_1 _09598_ (.A(_01767_),
    .B(_01768_),
    .Y(_01769_));
 sky130_fd_sc_hd__xnor2_1 _09599_ (.A(_01765_),
    .B(_01769_),
    .Y(_01770_));
 sky130_fd_sc_hd__nor3_1 _09600_ (.A(_01302_),
    .B(_01620_),
    .C(_01770_),
    .Y(_01771_));
 sky130_fd_sc_hd__o21a_1 _09601_ (.A1(_01302_),
    .A2(_01620_),
    .B1(_01770_),
    .X(_01772_));
 sky130_fd_sc_hd__or2_2 _09602_ (.A(_01771_),
    .B(_01772_),
    .X(_01773_));
 sky130_fd_sc_hd__a22oi_1 _09603_ (.A1(_06428_),
    .A2(_00415_),
    .B1(_00574_),
    .B2(_06439_),
    .Y(_01774_));
 sky130_fd_sc_hd__and4_1 _09604_ (.A(_06417_),
    .B(_00138_),
    .C(_00414_),
    .D(_00574_),
    .X(_01775_));
 sky130_fd_sc_hd__or2_1 _09605_ (.A(_01774_),
    .B(_01775_),
    .X(_01776_));
 sky130_fd_sc_hd__nand2_1 _09606_ (.A(_03059_),
    .B(_01600_),
    .Y(_01778_));
 sky130_fd_sc_hd__xnor2_1 _09607_ (.A(_01776_),
    .B(_01778_),
    .Y(_01779_));
 sky130_fd_sc_hd__clkbuf_4 _09608_ (.A(_01585_),
    .X(_01780_));
 sky130_fd_sc_hd__a32o_1 _09609_ (.A1(_02040_),
    .A2(_01600_),
    .A3(_01598_),
    .B1(_01597_),
    .B2(_00415_),
    .X(_01781_));
 sky130_fd_sc_hd__and3_1 _09610_ (.A(_02280_),
    .B(_01780_),
    .C(_01781_),
    .X(_01782_));
 sky130_fd_sc_hd__a21oi_1 _09611_ (.A1(_02335_),
    .A2(_01780_),
    .B1(_01781_),
    .Y(_01783_));
 sky130_fd_sc_hd__nor3_1 _09612_ (.A(_01779_),
    .B(_01782_),
    .C(_01783_),
    .Y(_01784_));
 sky130_fd_sc_hd__o21a_1 _09613_ (.A1(_01782_),
    .A2(_01783_),
    .B1(_01779_),
    .X(_01785_));
 sky130_fd_sc_hd__nor2_1 _09614_ (.A(_01784_),
    .B(_01785_),
    .Y(_01786_));
 sky130_fd_sc_hd__nand2_1 _09615_ (.A(_01605_),
    .B(_01786_),
    .Y(_01787_));
 sky130_fd_sc_hd__or2_1 _09616_ (.A(_01605_),
    .B(_01786_),
    .X(_01789_));
 sky130_fd_sc_hd__nand2_1 _09617_ (.A(_01787_),
    .B(_01789_),
    .Y(_01790_));
 sky130_fd_sc_hd__nand2_1 _09618_ (.A(_01582_),
    .B(_01594_),
    .Y(_01791_));
 sky130_fd_sc_hd__and3_1 _09619_ (.A(_01261_),
    .B(_01576_),
    .C(_01579_),
    .X(_01792_));
 sky130_fd_sc_hd__and3_1 _09620_ (.A(_01275_),
    .B(_01588_),
    .C(_01592_),
    .X(_01793_));
 sky130_fd_sc_hd__xnor2_1 _09621_ (.A(_01792_),
    .B(_01793_),
    .Y(_01794_));
 sky130_fd_sc_hd__xor2_1 _09622_ (.A(_01791_),
    .B(_01794_),
    .X(_01795_));
 sky130_fd_sc_hd__xnor2_1 _09623_ (.A(_01790_),
    .B(_01795_),
    .Y(_01796_));
 sky130_fd_sc_hd__or2_1 _09624_ (.A(_01573_),
    .B(_01595_),
    .X(_01797_));
 sky130_fd_sc_hd__and2_1 _09625_ (.A(_01573_),
    .B(_01595_),
    .X(_01798_));
 sky130_fd_sc_hd__a21o_1 _09626_ (.A1(_01797_),
    .A2(_01607_),
    .B1(_01798_),
    .X(_01800_));
 sky130_fd_sc_hd__and2b_1 _09627_ (.A_N(_01796_),
    .B(_01800_),
    .X(_01801_));
 sky130_fd_sc_hd__or2b_1 _09628_ (.A(_01800_),
    .B_N(_01796_),
    .X(_01802_));
 sky130_fd_sc_hd__and2b_1 _09629_ (.A_N(_01801_),
    .B(_01802_),
    .X(_01803_));
 sky130_fd_sc_hd__or2b_1 _09630_ (.A(_01608_),
    .B_N(_01609_),
    .X(_01804_));
 sky130_fd_sc_hd__a21bo_1 _09631_ (.A1(_01610_),
    .A2(_01612_),
    .B1_N(_01804_),
    .X(_01805_));
 sky130_fd_sc_hd__xnor2_2 _09632_ (.A(_01803_),
    .B(_01805_),
    .Y(_01806_));
 sky130_fd_sc_hd__xnor2_2 _09633_ (.A(_01773_),
    .B(_01806_),
    .Y(_01807_));
 sky130_fd_sc_hd__and3_1 _09634_ (.A(_01197_),
    .B(_04510_),
    .C(net18),
    .X(_01808_));
 sky130_fd_sc_hd__a22o_1 _09635_ (.A1(_01197_),
    .A2(_01177_),
    .B1(_01246_),
    .B2(_04510_),
    .X(_01809_));
 sky130_fd_sc_hd__a21bo_1 _09636_ (.A1(_01177_),
    .A2(_01808_),
    .B1_N(_01809_),
    .X(_01811_));
 sky130_fd_sc_hd__nand2_1 _09637_ (.A(_01744_),
    .B(net19),
    .Y(_01812_));
 sky130_fd_sc_hd__xor2_1 _09638_ (.A(_01811_),
    .B(_01812_),
    .X(_01813_));
 sky130_fd_sc_hd__a31o_1 _09639_ (.A1(_00300_),
    .A2(net19),
    .A3(_01565_),
    .B1(_01567_),
    .X(_01814_));
 sky130_fd_sc_hd__nand2_1 _09640_ (.A(_00311_),
    .B(net20),
    .Y(_01815_));
 sky130_fd_sc_hd__xnor2_1 _09641_ (.A(_01814_),
    .B(_01815_),
    .Y(_01816_));
 sky130_fd_sc_hd__xnor2_1 _09642_ (.A(_01813_),
    .B(_01816_),
    .Y(_01817_));
 sky130_fd_sc_hd__nor3_1 _09643_ (.A(_01255_),
    .B(_01571_),
    .C(_01817_),
    .Y(_01818_));
 sky130_fd_sc_hd__o21a_1 _09644_ (.A1(_01255_),
    .A2(_01571_),
    .B1(_01817_),
    .X(_01819_));
 sky130_fd_sc_hd__or2_2 _09645_ (.A(_01818_),
    .B(_01819_),
    .X(_01820_));
 sky130_fd_sc_hd__xnor2_4 _09646_ (.A(_01807_),
    .B(_01820_),
    .Y(_01822_));
 sky130_fd_sc_hd__o21a_1 _09647_ (.A1(_01614_),
    .A2(_01621_),
    .B1(_01572_),
    .X(_01823_));
 sky130_fd_sc_hd__a21o_2 _09648_ (.A1(_01614_),
    .A2(_01621_),
    .B1(_01823_),
    .X(_01824_));
 sky130_fd_sc_hd__xor2_4 _09649_ (.A(_01822_),
    .B(_01824_),
    .X(_01825_));
 sky130_fd_sc_hd__and2_1 _09650_ (.A(_01563_),
    .B(_01623_),
    .X(_01826_));
 sky130_fd_sc_hd__a21o_2 _09651_ (.A1(_01307_),
    .A2(_01625_),
    .B1(_01826_),
    .X(_01827_));
 sky130_fd_sc_hd__xor2_4 _09652_ (.A(_01825_),
    .B(_01827_),
    .X(_01828_));
 sky130_fd_sc_hd__or3b_2 _09653_ (.A(_01759_),
    .B(_01760_),
    .C_N(_01828_),
    .X(_01829_));
 sky130_fd_sc_hd__o21bai_2 _09654_ (.A1(_01759_),
    .A2(_01760_),
    .B1_N(_01828_),
    .Y(_01830_));
 sky130_fd_sc_hd__o21ba_1 _09655_ (.A1(_01626_),
    .A2(_01561_),
    .B1_N(_01560_),
    .X(_01831_));
 sky130_fd_sc_hd__nand3_4 _09656_ (.A(_01829_),
    .B(_01830_),
    .C(_01831_),
    .Y(_01833_));
 sky130_fd_sc_hd__a21o_1 _09657_ (.A1(_01829_),
    .A2(_01830_),
    .B1(_01831_),
    .X(_01834_));
 sky130_fd_sc_hd__nand3_1 _09658_ (.A(_01631_),
    .B(_01833_),
    .C(_01834_),
    .Y(_01835_));
 sky130_fd_sc_hd__a21o_1 _09659_ (.A1(_01833_),
    .A2(_01834_),
    .B1(_01631_),
    .X(_01836_));
 sky130_fd_sc_hd__and2_2 _09660_ (.A(_01835_),
    .B(_01836_),
    .X(_01837_));
 sky130_fd_sc_hd__xor2_4 _09661_ (.A(_01649_),
    .B(_01837_),
    .X(net84));
 sky130_fd_sc_hd__nor2_1 _09662_ (.A(_01740_),
    .B(_01741_),
    .Y(_01838_));
 sky130_fd_sc_hd__nand2_1 _09663_ (.A(_00670_),
    .B(_00145_),
    .Y(_01839_));
 sky130_fd_sc_hd__a21boi_1 _09664_ (.A1(_00843_),
    .A2(_00635_),
    .B1_N(_01839_),
    .Y(_01840_));
 sky130_fd_sc_hd__and4_1 _09665_ (.A(_00843_),
    .B(_00670_),
    .C(_00145_),
    .D(_04917_),
    .X(_01841_));
 sky130_fd_sc_hd__nor2_1 _09666_ (.A(_01840_),
    .B(_01841_),
    .Y(_01843_));
 sky130_fd_sc_hd__and3_1 _09667_ (.A(_00654_),
    .B(_00859_),
    .C(_01843_),
    .X(_01844_));
 sky130_fd_sc_hd__a21oi_1 _09668_ (.A1(_00654_),
    .A2(_00859_),
    .B1(_01843_),
    .Y(_01845_));
 sky130_fd_sc_hd__nor2_1 _09669_ (.A(_01844_),
    .B(_01845_),
    .Y(_01846_));
 sky130_fd_sc_hd__o21a_1 _09670_ (.A1(_01724_),
    .A2(_01726_),
    .B1(_01846_),
    .X(_01847_));
 sky130_fd_sc_hd__nor3_1 _09671_ (.A(_01724_),
    .B(_01726_),
    .C(_01846_),
    .Y(_01848_));
 sky130_fd_sc_hd__nor2_1 _09672_ (.A(_01847_),
    .B(_01848_),
    .Y(_01849_));
 sky130_fd_sc_hd__o21a_1 _09673_ (.A1(_01729_),
    .A2(net143),
    .B1(_01849_),
    .X(_01850_));
 sky130_fd_sc_hd__nor3_1 _09674_ (.A(_01729_),
    .B(net143),
    .C(_01849_),
    .Y(_01851_));
 sky130_fd_sc_hd__nor2_1 _09675_ (.A(_01850_),
    .B(_01851_),
    .Y(_01852_));
 sky130_fd_sc_hd__xnor2_1 _09676_ (.A(_01735_),
    .B(_01852_),
    .Y(_01854_));
 sky130_fd_sc_hd__and2_1 _09677_ (.A(_01838_),
    .B(_01854_),
    .X(_01855_));
 sky130_fd_sc_hd__nor2_1 _09678_ (.A(_01838_),
    .B(_01854_),
    .Y(_01856_));
 sky130_fd_sc_hd__nor2_1 _09679_ (.A(_01855_),
    .B(_01856_),
    .Y(_01857_));
 sky130_fd_sc_hd__o21a_1 _09680_ (.A1(_01737_),
    .A2(_01746_),
    .B1(_01743_),
    .X(_01858_));
 sky130_fd_sc_hd__and2_1 _09681_ (.A(_01857_),
    .B(_01858_),
    .X(_01859_));
 sky130_fd_sc_hd__nor2_1 _09682_ (.A(_01857_),
    .B(_01858_),
    .Y(_01860_));
 sky130_fd_sc_hd__nor2_1 _09683_ (.A(_01859_),
    .B(_01860_),
    .Y(_01861_));
 sky130_fd_sc_hd__inv_2 _09684_ (.A(_01861_),
    .Y(_01862_));
 sky130_fd_sc_hd__a31o_1 _09685_ (.A1(_01720_),
    .A2(_01485_),
    .A3(_01750_),
    .B1(_01749_),
    .X(_01863_));
 sky130_fd_sc_hd__nor2_1 _09686_ (.A(_01862_),
    .B(_01863_),
    .Y(_01865_));
 sky130_fd_sc_hd__and2_1 _09687_ (.A(_01862_),
    .B(_01863_),
    .X(_01866_));
 sky130_fd_sc_hd__nor2_2 _09688_ (.A(_01865_),
    .B(_01866_),
    .Y(_01867_));
 sky130_fd_sc_hd__xnor2_2 _09689_ (.A(_01754_),
    .B(_01867_),
    .Y(_01868_));
 sky130_fd_sc_hd__nand2_1 _09690_ (.A(_04939_),
    .B(_00379_),
    .Y(_01869_));
 sky130_fd_sc_hd__and3_1 _09691_ (.A(_05181_),
    .B(_04059_),
    .C(_01705_),
    .X(_01870_));
 sky130_fd_sc_hd__nor2_1 _09692_ (.A(_01703_),
    .B(_01707_),
    .Y(_01871_));
 sky130_fd_sc_hd__a31o_1 _09693_ (.A1(_05192_),
    .A2(_00373_),
    .A3(_01701_),
    .B1(_01699_),
    .X(_01872_));
 sky130_fd_sc_hd__a22oi_1 _09694_ (.A1(_04378_),
    .A2(_04103_),
    .B1(_00777_),
    .B2(_02971_),
    .Y(_01873_));
 sky130_fd_sc_hd__and4_1 _09695_ (.A(_02960_),
    .B(_04367_),
    .C(_04180_),
    .D(_04191_),
    .X(_01874_));
 sky130_fd_sc_hd__nor2_1 _09696_ (.A(_01873_),
    .B(_01874_),
    .Y(_01876_));
 sky130_fd_sc_hd__nand2_1 _09697_ (.A(_04598_),
    .B(_04026_),
    .Y(_01877_));
 sky130_fd_sc_hd__xnor2_1 _09698_ (.A(_01876_),
    .B(_01877_),
    .Y(_01878_));
 sky130_fd_sc_hd__xor2_1 _09699_ (.A(_01872_),
    .B(_01878_),
    .X(_01879_));
 sky130_fd_sc_hd__o21a_1 _09700_ (.A1(_01870_),
    .A2(_01871_),
    .B1(_01879_),
    .X(_01880_));
 sky130_fd_sc_hd__or3_1 _09701_ (.A(_01870_),
    .B(_01871_),
    .C(_01879_),
    .X(_01881_));
 sky130_fd_sc_hd__or2b_1 _09702_ (.A(_01880_),
    .B_N(_01881_),
    .X(_01882_));
 sky130_fd_sc_hd__xnor2_1 _09703_ (.A(_01709_),
    .B(_01882_),
    .Y(_01883_));
 sky130_fd_sc_hd__and2_1 _09704_ (.A(_00388_),
    .B(_00459_),
    .X(_01884_));
 sky130_fd_sc_hd__nand2_1 _09705_ (.A(_01883_),
    .B(_01884_),
    .Y(_01885_));
 sky130_fd_sc_hd__or2_1 _09706_ (.A(_01883_),
    .B(_01884_),
    .X(_01887_));
 sky130_fd_sc_hd__nand2_1 _09707_ (.A(_01885_),
    .B(_01887_),
    .Y(_01888_));
 sky130_fd_sc_hd__xor2_2 _09708_ (.A(_01869_),
    .B(_01888_),
    .X(_01889_));
 sky130_fd_sc_hd__nor2_1 _09709_ (.A(_01682_),
    .B(_01683_),
    .Y(_01890_));
 sky130_fd_sc_hd__o21ba_1 _09710_ (.A1(_01665_),
    .A2(_01669_),
    .B1_N(_01666_),
    .X(_01891_));
 sky130_fd_sc_hd__a22o_1 _09711_ (.A1(_06461_),
    .A2(_01508_),
    .B1(_01505_),
    .B2(_02160_),
    .X(_01892_));
 sky130_fd_sc_hd__and4_1 _09712_ (.A(_02160_),
    .B(_06461_),
    .C(_01508_),
    .D(_01504_),
    .X(_01893_));
 sky130_fd_sc_hd__inv_2 _09713_ (.A(_01893_),
    .Y(_01894_));
 sky130_fd_sc_hd__a22oi_1 _09714_ (.A1(_06494_),
    .A2(_00608_),
    .B1(_01892_),
    .B2(_01894_),
    .Y(_01895_));
 sky130_fd_sc_hd__and4_1 _09715_ (.A(_06483_),
    .B(_00607_),
    .C(_01892_),
    .D(_01894_),
    .X(_01896_));
 sky130_fd_sc_hd__nor2_1 _09716_ (.A(_01895_),
    .B(_01896_),
    .Y(_01898_));
 sky130_fd_sc_hd__xnor2_1 _09717_ (.A(_01891_),
    .B(_01898_),
    .Y(_01899_));
 sky130_fd_sc_hd__o21a_1 _09718_ (.A1(_01672_),
    .A2(_01674_),
    .B1(_01899_),
    .X(_01900_));
 sky130_fd_sc_hd__nor3_1 _09719_ (.A(_01672_),
    .B(_01674_),
    .C(_01899_),
    .Y(_01901_));
 sky130_fd_sc_hd__nor2_1 _09720_ (.A(_01900_),
    .B(_01901_),
    .Y(_01902_));
 sky130_fd_sc_hd__xnor2_1 _09721_ (.A(_01677_),
    .B(_01902_),
    .Y(_01903_));
 sky130_fd_sc_hd__and2_1 _09722_ (.A(_01890_),
    .B(_01903_),
    .X(_01904_));
 sky130_fd_sc_hd__nor2_1 _09723_ (.A(_01890_),
    .B(_01903_),
    .Y(_01905_));
 sky130_fd_sc_hd__or2_1 _09724_ (.A(_01904_),
    .B(_01905_),
    .X(_01906_));
 sky130_fd_sc_hd__o21a_1 _09725_ (.A1(_01681_),
    .A2(_01684_),
    .B1(_01680_),
    .X(_01907_));
 sky130_fd_sc_hd__a21o_1 _09726_ (.A1(_01681_),
    .A2(_01684_),
    .B1(_01907_),
    .X(_01909_));
 sky130_fd_sc_hd__nor2_1 _09727_ (.A(_01906_),
    .B(_01909_),
    .Y(_01910_));
 sky130_fd_sc_hd__and2_1 _09728_ (.A(_01906_),
    .B(_01909_),
    .X(_01911_));
 sky130_fd_sc_hd__nor2_2 _09729_ (.A(_01910_),
    .B(_01911_),
    .Y(_01912_));
 sky130_fd_sc_hd__or2b_1 _09730_ (.A(_01686_),
    .B_N(_01688_),
    .X(_01913_));
 sky130_fd_sc_hd__a31o_1 _09731_ (.A1(_01539_),
    .A2(_01693_),
    .A3(_01913_),
    .B1(_01691_),
    .X(_01914_));
 sky130_fd_sc_hd__a31o_2 _09732_ (.A1(_01541_),
    .A2(_01543_),
    .A3(_01692_),
    .B1(_01914_),
    .X(_01915_));
 sky130_fd_sc_hd__xor2_2 _09733_ (.A(_01912_),
    .B(_01915_),
    .X(_01916_));
 sky130_fd_sc_hd__nand2_1 _09734_ (.A(_02467_),
    .B(_01060_),
    .Y(_01917_));
 sky130_fd_sc_hd__and3_1 _09735_ (.A(_01339_),
    .B(_01058_),
    .C(_01657_),
    .X(_01918_));
 sky130_fd_sc_hd__nor2_1 _09736_ (.A(_01654_),
    .B(_01659_),
    .Y(_01920_));
 sky130_fd_sc_hd__a31o_1 _09737_ (.A1(_04081_),
    .A2(_01410_),
    .A3(_01652_),
    .B1(_01651_),
    .X(_01921_));
 sky130_fd_sc_hd__a22oi_1 _09738_ (.A1(_00891_),
    .A2(_01545_),
    .B1(net52),
    .B2(_03587_),
    .Y(_01922_));
 sky130_fd_sc_hd__and4_1 _09739_ (.A(_04169_),
    .B(_01076_),
    .C(_01545_),
    .D(net52),
    .X(_01923_));
 sky130_fd_sc_hd__nor2_1 _09740_ (.A(_01922_),
    .B(_01923_),
    .Y(_01924_));
 sky130_fd_sc_hd__nand2_1 _09741_ (.A(_04268_),
    .B(net50),
    .Y(_01925_));
 sky130_fd_sc_hd__xnor2_1 _09742_ (.A(_01924_),
    .B(_01925_),
    .Y(_01926_));
 sky130_fd_sc_hd__xor2_1 _09743_ (.A(_01921_),
    .B(_01926_),
    .X(_01927_));
 sky130_fd_sc_hd__o21a_1 _09744_ (.A1(_01918_),
    .A2(_01920_),
    .B1(_01927_),
    .X(_01928_));
 sky130_fd_sc_hd__or3_1 _09745_ (.A(_01918_),
    .B(_01920_),
    .C(_01927_),
    .X(_01929_));
 sky130_fd_sc_hd__or2b_1 _09746_ (.A(_01928_),
    .B_N(_01929_),
    .X(_01931_));
 sky130_fd_sc_hd__xnor2_1 _09747_ (.A(_01661_),
    .B(_01931_),
    .Y(_01932_));
 sky130_fd_sc_hd__clkbuf_4 _09748_ (.A(net53),
    .X(_01933_));
 sky130_fd_sc_hd__clkbuf_4 _09749_ (.A(_01933_),
    .X(_01934_));
 sky130_fd_sc_hd__and2_1 _09750_ (.A(_00453_),
    .B(_01934_),
    .X(_01935_));
 sky130_fd_sc_hd__nand2_1 _09751_ (.A(_01932_),
    .B(_01935_),
    .Y(_01936_));
 sky130_fd_sc_hd__or2_1 _09752_ (.A(_01932_),
    .B(_01935_),
    .X(_01937_));
 sky130_fd_sc_hd__nand2_1 _09753_ (.A(_01936_),
    .B(_01937_),
    .Y(_01938_));
 sky130_fd_sc_hd__xor2_2 _09754_ (.A(_01917_),
    .B(_01938_),
    .X(_01939_));
 sky130_fd_sc_hd__xor2_1 _09755_ (.A(_01916_),
    .B(_01939_),
    .X(_01940_));
 sky130_fd_sc_hd__xnor2_1 _09756_ (.A(_01889_),
    .B(_01940_),
    .Y(_01942_));
 sky130_fd_sc_hd__o21a_1 _09757_ (.A1(_01663_),
    .A2(_01696_),
    .B1(_01712_),
    .X(_01943_));
 sky130_fd_sc_hd__a21o_1 _09758_ (.A1(_01663_),
    .A2(_01696_),
    .B1(_01943_),
    .X(_01944_));
 sky130_fd_sc_hd__xor2_1 _09759_ (.A(_01942_),
    .B(_01944_),
    .X(_01945_));
 sky130_fd_sc_hd__nor2_1 _09760_ (.A(_01713_),
    .B(_01715_),
    .Y(_01946_));
 sky130_fd_sc_hd__a211oi_1 _09761_ (.A1(_01716_),
    .A2(_01717_),
    .B1(_01945_),
    .C1(_01946_),
    .Y(_01947_));
 sky130_fd_sc_hd__and2_2 _09762_ (.A(_01946_),
    .B(_01945_),
    .X(_01948_));
 sky130_fd_sc_hd__and3_2 _09763_ (.A(_01716_),
    .B(_01717_),
    .C(_01945_),
    .X(_01949_));
 sky130_fd_sc_hd__nor3_2 _09764_ (.A(_01947_),
    .B(_01948_),
    .C(_01949_),
    .Y(_01950_));
 sky130_fd_sc_hd__xor2_2 _09765_ (.A(_01868_),
    .B(_01950_),
    .X(_01951_));
 sky130_fd_sc_hd__buf_2 _09766_ (.A(net21),
    .X(_01953_));
 sky130_fd_sc_hd__clkbuf_4 _09767_ (.A(_01953_),
    .X(_01954_));
 sky130_fd_sc_hd__buf_4 _09768_ (.A(_01954_),
    .X(_01955_));
 sky130_fd_sc_hd__clkbuf_4 _09769_ (.A(_01955_),
    .X(_01956_));
 sky130_fd_sc_hd__clkbuf_4 _09770_ (.A(_01956_),
    .X(_01957_));
 sky130_fd_sc_hd__buf_4 _09771_ (.A(_01957_),
    .X(_01958_));
 sky130_fd_sc_hd__nand2_1 _09772_ (.A(_00344_),
    .B(_01958_),
    .Y(_01959_));
 sky130_fd_sc_hd__clkbuf_4 _09773_ (.A(net20),
    .X(_01960_));
 sky130_fd_sc_hd__and3_1 _09774_ (.A(_00322_),
    .B(_01960_),
    .C(_01814_),
    .X(_01961_));
 sky130_fd_sc_hd__and2_1 _09775_ (.A(_01813_),
    .B(_01816_),
    .X(_01962_));
 sky130_fd_sc_hd__o2bb2ai_1 _09776_ (.A1_N(_01178_),
    .A2_N(_01808_),
    .B1(_01811_),
    .B2(_01812_),
    .Y(_01964_));
 sky130_fd_sc_hd__nand2_1 _09777_ (.A(_01295_),
    .B(_01246_),
    .Y(_01965_));
 sky130_fd_sc_hd__nand2_1 _09778_ (.A(_01306_),
    .B(net19),
    .Y(_01966_));
 sky130_fd_sc_hd__and4_1 _09779_ (.A(_01197_),
    .B(_04510_),
    .C(_01246_),
    .D(net19),
    .X(_01967_));
 sky130_fd_sc_hd__a21oi_1 _09780_ (.A1(_01965_),
    .A2(_01966_),
    .B1(_01967_),
    .Y(_01968_));
 sky130_fd_sc_hd__nand2_1 _09781_ (.A(_01744_),
    .B(net20),
    .Y(_01969_));
 sky130_fd_sc_hd__xnor2_1 _09782_ (.A(_01968_),
    .B(_01969_),
    .Y(_01970_));
 sky130_fd_sc_hd__xor2_1 _09783_ (.A(_01964_),
    .B(_01970_),
    .X(_01971_));
 sky130_fd_sc_hd__o21a_1 _09784_ (.A1(_01961_),
    .A2(_01962_),
    .B1(_01971_),
    .X(_01972_));
 sky130_fd_sc_hd__or3_1 _09785_ (.A(_01961_),
    .B(_01962_),
    .C(_01971_),
    .X(_01973_));
 sky130_fd_sc_hd__and2b_1 _09786_ (.A_N(_01972_),
    .B(_01973_),
    .X(_01975_));
 sky130_fd_sc_hd__xor2_1 _09787_ (.A(_01818_),
    .B(_01975_),
    .X(_01976_));
 sky130_fd_sc_hd__and3_1 _09788_ (.A(_02456_),
    .B(_01180_),
    .C(_01976_),
    .X(_01977_));
 sky130_fd_sc_hd__a21o_1 _09789_ (.A1(_02456_),
    .A2(_01181_),
    .B1(_01976_),
    .X(_01978_));
 sky130_fd_sc_hd__and2b_1 _09790_ (.A_N(_01977_),
    .B(_01978_),
    .X(_01979_));
 sky130_fd_sc_hd__xnor2_2 _09791_ (.A(_01959_),
    .B(_01979_),
    .Y(_01980_));
 sky130_fd_sc_hd__nor2_1 _09792_ (.A(_01792_),
    .B(_01793_),
    .Y(_01981_));
 sky130_fd_sc_hd__o21ba_1 _09793_ (.A1(_01774_),
    .A2(_01778_),
    .B1_N(_01775_),
    .X(_01982_));
 sky130_fd_sc_hd__a22o_1 _09794_ (.A1(_06417_),
    .A2(_00574_),
    .B1(_01600_),
    .B2(_06439_),
    .X(_01983_));
 sky130_fd_sc_hd__and4_1 _09795_ (.A(_05456_),
    .B(_00138_),
    .C(_00572_),
    .D(_01586_),
    .X(_01984_));
 sky130_fd_sc_hd__inv_2 _09796_ (.A(_01984_),
    .Y(_01986_));
 sky130_fd_sc_hd__a22oi_1 _09797_ (.A1(_03070_),
    .A2(_01585_),
    .B1(_01983_),
    .B2(_01986_),
    .Y(_01987_));
 sky130_fd_sc_hd__and4_1 _09798_ (.A(_03059_),
    .B(_01585_),
    .C(_01983_),
    .D(_01986_),
    .X(_01988_));
 sky130_fd_sc_hd__nor2_1 _09799_ (.A(_01987_),
    .B(_01988_),
    .Y(_01989_));
 sky130_fd_sc_hd__xnor2_1 _09800_ (.A(_01982_),
    .B(_01989_),
    .Y(_01990_));
 sky130_fd_sc_hd__o21a_1 _09801_ (.A1(_01782_),
    .A2(_01784_),
    .B1(_01990_),
    .X(_01991_));
 sky130_fd_sc_hd__nor3_1 _09802_ (.A(_01782_),
    .B(_01784_),
    .C(_01990_),
    .Y(_01992_));
 sky130_fd_sc_hd__nor2_1 _09803_ (.A(_01991_),
    .B(_01992_),
    .Y(_01993_));
 sky130_fd_sc_hd__xnor2_1 _09804_ (.A(_01787_),
    .B(_01993_),
    .Y(_01994_));
 sky130_fd_sc_hd__and2_1 _09805_ (.A(_01981_),
    .B(_01994_),
    .X(_01995_));
 sky130_fd_sc_hd__nor2_1 _09806_ (.A(_01981_),
    .B(_01994_),
    .Y(_01997_));
 sky130_fd_sc_hd__or2_1 _09807_ (.A(_01995_),
    .B(_01997_),
    .X(_01998_));
 sky130_fd_sc_hd__o21a_1 _09808_ (.A1(_01791_),
    .A2(_01794_),
    .B1(_01790_),
    .X(_01999_));
 sky130_fd_sc_hd__a21o_1 _09809_ (.A1(_01791_),
    .A2(_01794_),
    .B1(_01999_),
    .X(_02000_));
 sky130_fd_sc_hd__nor2_1 _09810_ (.A(_01998_),
    .B(_02000_),
    .Y(_02001_));
 sky130_fd_sc_hd__and2_1 _09811_ (.A(_01998_),
    .B(_02000_),
    .X(_02002_));
 sky130_fd_sc_hd__nor2_2 _09812_ (.A(_02001_),
    .B(_02002_),
    .Y(_02003_));
 sky130_fd_sc_hd__o21ai_1 _09813_ (.A1(_01804_),
    .A2(_01801_),
    .B1(_01802_),
    .Y(_02004_));
 sky130_fd_sc_hd__a31o_4 _09814_ (.A1(_01610_),
    .A2(_01612_),
    .A3(_01803_),
    .B1(_02004_),
    .X(_02005_));
 sky130_fd_sc_hd__xor2_2 _09815_ (.A(_02003_),
    .B(_02005_),
    .X(_02006_));
 sky130_fd_sc_hd__buf_4 _09816_ (.A(_01188_),
    .X(_02008_));
 sky130_fd_sc_hd__nand2_1 _09817_ (.A(_00530_),
    .B(_02008_),
    .Y(_02009_));
 sky130_fd_sc_hd__and3_1 _09818_ (.A(_00486_),
    .B(_01260_),
    .C(_01767_),
    .X(_02010_));
 sky130_fd_sc_hd__and2_1 _09819_ (.A(_01765_),
    .B(_01769_),
    .X(_02011_));
 sky130_fd_sc_hd__o2bb2ai_1 _09820_ (.A1_N(_03696_),
    .A2_N(_01761_),
    .B1(_01763_),
    .B2(_01764_),
    .Y(_02012_));
 sky130_fd_sc_hd__nand2_1 _09821_ (.A(_06819_),
    .B(_00423_),
    .Y(_02013_));
 sky130_fd_sc_hd__nand2_1 _09822_ (.A(_06821_),
    .B(net10),
    .Y(_02014_));
 sky130_fd_sc_hd__and4_1 _09823_ (.A(_06818_),
    .B(_06820_),
    .C(net9),
    .D(net10),
    .X(_02015_));
 sky130_fd_sc_hd__a21oi_1 _09824_ (.A1(_02013_),
    .A2(_02014_),
    .B1(_02015_),
    .Y(_02016_));
 sky130_fd_sc_hd__nand2_1 _09825_ (.A(_03510_),
    .B(net11),
    .Y(_02017_));
 sky130_fd_sc_hd__xnor2_1 _09826_ (.A(_02016_),
    .B(_02017_),
    .Y(_02019_));
 sky130_fd_sc_hd__xor2_1 _09827_ (.A(_02012_),
    .B(_02019_),
    .X(_02020_));
 sky130_fd_sc_hd__o21a_1 _09828_ (.A1(_02010_),
    .A2(_02011_),
    .B1(_02020_),
    .X(_02021_));
 sky130_fd_sc_hd__or3_1 _09829_ (.A(_02010_),
    .B(_02011_),
    .C(_02020_),
    .X(_02022_));
 sky130_fd_sc_hd__and2b_1 _09830_ (.A_N(_02021_),
    .B(_02022_),
    .X(_02023_));
 sky130_fd_sc_hd__xor2_1 _09831_ (.A(_01771_),
    .B(_02023_),
    .X(_02024_));
 sky130_fd_sc_hd__and3_1 _09832_ (.A(_07004_),
    .B(_00390_),
    .C(_02024_),
    .X(_02025_));
 sky130_fd_sc_hd__a21o_1 _09833_ (.A1(_07004_),
    .A2(_00390_),
    .B1(_02024_),
    .X(_02026_));
 sky130_fd_sc_hd__and2b_1 _09834_ (.A_N(_02025_),
    .B(_02026_),
    .X(_02027_));
 sky130_fd_sc_hd__xnor2_2 _09835_ (.A(_02009_),
    .B(_02027_),
    .Y(_02028_));
 sky130_fd_sc_hd__xor2_1 _09836_ (.A(_02006_),
    .B(_02028_),
    .X(_02030_));
 sky130_fd_sc_hd__xnor2_2 _09837_ (.A(_01980_),
    .B(_02030_),
    .Y(_02031_));
 sky130_fd_sc_hd__o21a_1 _09838_ (.A1(_01773_),
    .A2(_01806_),
    .B1(_01820_),
    .X(_02032_));
 sky130_fd_sc_hd__a21o_1 _09839_ (.A1(_01773_),
    .A2(_01806_),
    .B1(_02032_),
    .X(_02033_));
 sky130_fd_sc_hd__xor2_1 _09840_ (.A(_02031_),
    .B(_02033_),
    .X(_02034_));
 sky130_fd_sc_hd__nor2_1 _09841_ (.A(_01822_),
    .B(_01824_),
    .Y(_02035_));
 sky130_fd_sc_hd__a211oi_1 _09842_ (.A1(_01825_),
    .A2(_01827_),
    .B1(_02034_),
    .C1(_02035_),
    .Y(_02036_));
 sky130_fd_sc_hd__and2_2 _09843_ (.A(_02035_),
    .B(_02034_),
    .X(_02037_));
 sky130_fd_sc_hd__and3_2 _09844_ (.A(_01825_),
    .B(_01827_),
    .C(_02034_),
    .X(_02038_));
 sky130_fd_sc_hd__or3_4 _09845_ (.A(_02036_),
    .B(_02037_),
    .C(_02038_),
    .X(_02039_));
 sky130_fd_sc_hd__xnor2_4 _09846_ (.A(_01951_),
    .B(_02039_),
    .Y(_02041_));
 sky130_fd_sc_hd__or2_1 _09847_ (.A(_01828_),
    .B(_01759_),
    .X(_02042_));
 sky130_fd_sc_hd__or2b_2 _09848_ (.A(_01760_),
    .B_N(_02042_),
    .X(_02043_));
 sky130_fd_sc_hd__xor2_4 _09849_ (.A(_02041_),
    .B(_02043_),
    .X(_02044_));
 sky130_fd_sc_hd__xor2_4 _09850_ (.A(_01833_),
    .B(_02044_),
    .X(_02045_));
 sky130_fd_sc_hd__and4_2 _09851_ (.A(_01633_),
    .B(_01634_),
    .C(_01835_),
    .D(_01836_),
    .X(_02046_));
 sky130_fd_sc_hd__o211ai_1 _09852_ (.A1(_01627_),
    .A2(_01628_),
    .B1(_01629_),
    .C1(_01630_),
    .Y(_02047_));
 sky130_fd_sc_hd__nand2_1 _09853_ (.A(_01833_),
    .B(_01834_),
    .Y(_02048_));
 sky130_fd_sc_hd__a21oi_4 _09854_ (.A1(_02047_),
    .A2(_01633_),
    .B1(_02048_),
    .Y(_02049_));
 sky130_fd_sc_hd__a21oi_1 _09855_ (.A1(_01640_),
    .A2(_02046_),
    .B1(_02049_),
    .Y(_02050_));
 sky130_fd_sc_hd__xnor2_1 _09856_ (.A(_02045_),
    .B(_02050_),
    .Y(net85));
 sky130_fd_sc_hd__and3b_2 _09857_ (.A_N(_01760_),
    .B(_02041_),
    .C(_02042_),
    .X(_02052_));
 sky130_fd_sc_hd__nand2_1 _09858_ (.A(_01868_),
    .B(_01950_),
    .Y(_02053_));
 sky130_fd_sc_hd__nor2_1 _09859_ (.A(_01868_),
    .B(_01950_),
    .Y(_02054_));
 sky130_fd_sc_hd__a21o_2 _09860_ (.A1(_02053_),
    .A2(_02039_),
    .B1(_02054_),
    .X(_02055_));
 sky130_fd_sc_hd__nor2_1 _09861_ (.A(_02031_),
    .B(_02033_),
    .Y(_02056_));
 sky130_fd_sc_hd__a21o_1 _09862_ (.A1(_00519_),
    .A2(_01188_),
    .B1(_02025_),
    .X(_02057_));
 sky130_fd_sc_hd__nand2_1 _09863_ (.A(_02026_),
    .B(_02057_),
    .Y(_02058_));
 sky130_fd_sc_hd__a22o_1 _09864_ (.A1(_00004_),
    .A2(_00390_),
    .B1(_00393_),
    .B2(_07004_),
    .X(_02059_));
 sky130_fd_sc_hd__nand4_2 _09865_ (.A(_06765_),
    .B(_06775_),
    .C(_03707_),
    .D(_03740_),
    .Y(_02060_));
 sky130_fd_sc_hd__nand2_1 _09866_ (.A(_02012_),
    .B(_02019_),
    .Y(_02062_));
 sky130_fd_sc_hd__a31o_1 _09867_ (.A1(_03521_),
    .A2(_01260_),
    .A3(_02016_),
    .B1(_02015_),
    .X(_02063_));
 sky130_fd_sc_hd__a22o_1 _09868_ (.A1(_06873_),
    .A2(_00755_),
    .B1(_01260_),
    .B2(_06875_),
    .X(_02064_));
 sky130_fd_sc_hd__nand4_2 _09869_ (.A(_06964_),
    .B(_00121_),
    .C(_00755_),
    .D(_00741_),
    .Y(_02065_));
 sky130_fd_sc_hd__nand2_1 _09870_ (.A(_02064_),
    .B(_02065_),
    .Y(_02066_));
 sky130_fd_sc_hd__xor2_1 _09871_ (.A(_02063_),
    .B(_02066_),
    .X(_02067_));
 sky130_fd_sc_hd__nor2_1 _09872_ (.A(_02062_),
    .B(_02067_),
    .Y(_02068_));
 sky130_fd_sc_hd__nand2_1 _09873_ (.A(_02062_),
    .B(_02067_),
    .Y(_02069_));
 sky130_fd_sc_hd__or2b_1 _09874_ (.A(_02068_),
    .B_N(_02069_),
    .X(_02070_));
 sky130_fd_sc_hd__a21o_1 _09875_ (.A1(_01771_),
    .A2(_02022_),
    .B1(_02021_),
    .X(_02071_));
 sky130_fd_sc_hd__xnor2_1 _09876_ (.A(_02070_),
    .B(_02071_),
    .Y(_02073_));
 sky130_fd_sc_hd__a21o_1 _09877_ (.A1(_02059_),
    .A2(_02060_),
    .B1(_02073_),
    .X(_02074_));
 sky130_fd_sc_hd__nand3_1 _09878_ (.A(_02073_),
    .B(_02059_),
    .C(_02060_),
    .Y(_02075_));
 sky130_fd_sc_hd__nand2_1 _09879_ (.A(_02074_),
    .B(_02075_),
    .Y(_02076_));
 sky130_fd_sc_hd__a22o_1 _09880_ (.A1(_03554_),
    .A2(_00416_),
    .B1(_01288_),
    .B2(_00508_),
    .X(_02077_));
 sky130_fd_sc_hd__and4_1 _09881_ (.A(_03521_),
    .B(_00486_),
    .C(_00413_),
    .D(_00572_),
    .X(_02078_));
 sky130_fd_sc_hd__inv_2 _09882_ (.A(_02078_),
    .Y(_02079_));
 sky130_fd_sc_hd__and2_1 _09883_ (.A(_02077_),
    .B(_02079_),
    .X(_02080_));
 sky130_fd_sc_hd__xor2_1 _09884_ (.A(_02076_),
    .B(_02080_),
    .X(_02081_));
 sky130_fd_sc_hd__nor2_1 _09885_ (.A(_02058_),
    .B(_02081_),
    .Y(_02082_));
 sky130_fd_sc_hd__and2_1 _09886_ (.A(_02058_),
    .B(_02081_),
    .X(_02084_));
 sky130_fd_sc_hd__or2_1 _09887_ (.A(_02082_),
    .B(_02084_),
    .X(_02085_));
 sky130_fd_sc_hd__inv_2 _09888_ (.A(_02085_),
    .Y(_02086_));
 sky130_fd_sc_hd__or2b_1 _09889_ (.A(_01982_),
    .B_N(_01989_),
    .X(_02087_));
 sky130_fd_sc_hd__clkbuf_4 _09890_ (.A(_01780_),
    .X(_02088_));
 sky130_fd_sc_hd__a31o_1 _09891_ (.A1(_03070_),
    .A2(_02088_),
    .A3(_01983_),
    .B1(_01984_),
    .X(_02089_));
 sky130_fd_sc_hd__clkbuf_4 _09892_ (.A(_01601_),
    .X(_02090_));
 sky130_fd_sc_hd__a22oi_1 _09893_ (.A1(_06626_),
    .A2(_02090_),
    .B1(_02088_),
    .B2(_06450_),
    .Y(_02091_));
 sky130_fd_sc_hd__and4_1 _09894_ (.A(_06626_),
    .B(_06450_),
    .C(_02090_),
    .D(_02088_),
    .X(_02092_));
 sky130_fd_sc_hd__nor2_1 _09895_ (.A(_02091_),
    .B(_02092_),
    .Y(_02093_));
 sky130_fd_sc_hd__and2_1 _09896_ (.A(_02089_),
    .B(_02093_),
    .X(_02095_));
 sky130_fd_sc_hd__nor2_1 _09897_ (.A(_02089_),
    .B(_02093_),
    .Y(_02096_));
 sky130_fd_sc_hd__nor2_1 _09898_ (.A(_02095_),
    .B(_02096_),
    .Y(_02097_));
 sky130_fd_sc_hd__xnor2_1 _09899_ (.A(_02087_),
    .B(_02097_),
    .Y(_02098_));
 sky130_fd_sc_hd__a31o_1 _09900_ (.A1(_01605_),
    .A2(_01786_),
    .A3(_01993_),
    .B1(_01991_),
    .X(_02099_));
 sky130_fd_sc_hd__nor2_1 _09901_ (.A(_02098_),
    .B(_02099_),
    .Y(_02100_));
 sky130_fd_sc_hd__and2_1 _09902_ (.A(_02098_),
    .B(_02099_),
    .X(_02101_));
 sky130_fd_sc_hd__nor2_1 _09903_ (.A(_02100_),
    .B(_02101_),
    .Y(_02102_));
 sky130_fd_sc_hd__or2_1 _09904_ (.A(_01995_),
    .B(_02102_),
    .X(_02103_));
 sky130_fd_sc_hd__nand2_1 _09905_ (.A(_01995_),
    .B(_02102_),
    .Y(_02104_));
 sky130_fd_sc_hd__nand2_1 _09906_ (.A(_02103_),
    .B(_02104_),
    .Y(_02106_));
 sky130_fd_sc_hd__a21o_1 _09907_ (.A1(_02003_),
    .A2(_02005_),
    .B1(_02001_),
    .X(_02107_));
 sky130_fd_sc_hd__xnor2_2 _09908_ (.A(_02106_),
    .B(_02107_),
    .Y(_02108_));
 sky130_fd_sc_hd__xnor2_1 _09909_ (.A(_02086_),
    .B(_02108_),
    .Y(_02109_));
 sky130_fd_sc_hd__a21o_1 _09910_ (.A1(_00333_),
    .A2(_01955_),
    .B1(_01977_),
    .X(_02110_));
 sky130_fd_sc_hd__nand2_1 _09911_ (.A(_01978_),
    .B(_02110_),
    .Y(_02111_));
 sky130_fd_sc_hd__a22o_1 _09912_ (.A1(_03070_),
    .A2(_01180_),
    .B1(_01249_),
    .B2(_02335_),
    .X(_02112_));
 sky130_fd_sc_hd__nand4_2 _09913_ (.A(_02007_),
    .B(_02040_),
    .C(_01179_),
    .D(_01254_),
    .Y(_02113_));
 sky130_fd_sc_hd__nand2_1 _09914_ (.A(_01964_),
    .B(_01970_),
    .Y(_02114_));
 sky130_fd_sc_hd__a31o_1 _09915_ (.A1(_02138_),
    .A2(_01960_),
    .A3(_01968_),
    .B1(_01967_),
    .X(_02115_));
 sky130_fd_sc_hd__clkbuf_4 _09916_ (.A(_01564_),
    .X(_02117_));
 sky130_fd_sc_hd__a22o_1 _09917_ (.A1(_01361_),
    .A2(_02117_),
    .B1(_01960_),
    .B2(_00159_),
    .X(_02118_));
 sky130_fd_sc_hd__clkbuf_4 _09918_ (.A(_02117_),
    .X(_02119_));
 sky130_fd_sc_hd__clkbuf_4 _09919_ (.A(_01960_),
    .X(_02120_));
 sky130_fd_sc_hd__nand4_2 _09920_ (.A(_01361_),
    .B(_00159_),
    .C(_02119_),
    .D(_02120_),
    .Y(_02121_));
 sky130_fd_sc_hd__nand2_1 _09921_ (.A(_02118_),
    .B(_02121_),
    .Y(_02122_));
 sky130_fd_sc_hd__xor2_1 _09922_ (.A(_02115_),
    .B(_02122_),
    .X(_02123_));
 sky130_fd_sc_hd__nor2_1 _09923_ (.A(_02114_),
    .B(_02123_),
    .Y(_02124_));
 sky130_fd_sc_hd__nand2_1 _09924_ (.A(_02114_),
    .B(_02123_),
    .Y(_02125_));
 sky130_fd_sc_hd__or2b_1 _09925_ (.A(_02124_),
    .B_N(_02125_),
    .X(_02126_));
 sky130_fd_sc_hd__a21o_1 _09926_ (.A1(_01818_),
    .A2(_01973_),
    .B1(_01972_),
    .X(_02128_));
 sky130_fd_sc_hd__xnor2_1 _09927_ (.A(_02126_),
    .B(_02128_),
    .Y(_02129_));
 sky130_fd_sc_hd__a21o_1 _09928_ (.A1(_02112_),
    .A2(_02113_),
    .B1(_02129_),
    .X(_02130_));
 sky130_fd_sc_hd__nand3_1 _09929_ (.A(_02129_),
    .B(_02112_),
    .C(_02113_),
    .Y(_02131_));
 sky130_fd_sc_hd__nand2_1 _09930_ (.A(_02130_),
    .B(_02131_),
    .Y(_02132_));
 sky130_fd_sc_hd__clkbuf_4 _09931_ (.A(net22),
    .X(_02133_));
 sky130_fd_sc_hd__buf_2 _09932_ (.A(_02133_),
    .X(_02134_));
 sky130_fd_sc_hd__clkbuf_4 _09933_ (.A(_02134_),
    .X(_02135_));
 sky130_fd_sc_hd__a22o_1 _09934_ (.A1(_02138_),
    .A2(_01954_),
    .B1(_02135_),
    .B2(_00333_),
    .X(_02136_));
 sky130_fd_sc_hd__and4_1 _09935_ (.A(_02127_),
    .B(_00322_),
    .C(net21),
    .D(_02133_),
    .X(_02137_));
 sky130_fd_sc_hd__inv_2 _09936_ (.A(_02137_),
    .Y(_02139_));
 sky130_fd_sc_hd__and2_1 _09937_ (.A(_02136_),
    .B(_02139_),
    .X(_02140_));
 sky130_fd_sc_hd__xor2_1 _09938_ (.A(_02132_),
    .B(_02140_),
    .X(_02141_));
 sky130_fd_sc_hd__nor2_1 _09939_ (.A(_02111_),
    .B(_02141_),
    .Y(_02142_));
 sky130_fd_sc_hd__and2_1 _09940_ (.A(_02111_),
    .B(_02141_),
    .X(_02143_));
 sky130_fd_sc_hd__or2_1 _09941_ (.A(_02142_),
    .B(_02143_),
    .X(_02144_));
 sky130_fd_sc_hd__xnor2_2 _09942_ (.A(_02109_),
    .B(_02144_),
    .Y(_02145_));
 sky130_fd_sc_hd__a21o_1 _09943_ (.A1(_02006_),
    .A2(_02028_),
    .B1(_01980_),
    .X(_02146_));
 sky130_fd_sc_hd__o21a_1 _09944_ (.A1(_02006_),
    .A2(_02028_),
    .B1(_02146_),
    .X(_02147_));
 sky130_fd_sc_hd__xnor2_2 _09945_ (.A(_02145_),
    .B(_02147_),
    .Y(_02148_));
 sky130_fd_sc_hd__o31ai_4 _09946_ (.A1(_02056_),
    .A2(_02037_),
    .A3(_02038_),
    .B1(_02148_),
    .Y(_02150_));
 sky130_fd_sc_hd__o41a_4 _09947_ (.A1(_02056_),
    .A2(_02037_),
    .A3(_02038_),
    .A4(_02148_),
    .B1(_02150_),
    .X(_02151_));
 sky130_fd_sc_hd__nor2_1 _09948_ (.A(_01942_),
    .B(_01944_),
    .Y(_02152_));
 sky130_fd_sc_hd__a21bo_1 _09949_ (.A1(_01917_),
    .A2(_01936_),
    .B1_N(_01937_),
    .X(_02153_));
 sky130_fd_sc_hd__nand2_1 _09950_ (.A(_01921_),
    .B(_01926_),
    .Y(_02154_));
 sky130_fd_sc_hd__a31o_1 _09951_ (.A1(_01339_),
    .A2(_01410_),
    .A3(_01924_),
    .B1(_01923_),
    .X(_02155_));
 sky130_fd_sc_hd__buf_2 _09952_ (.A(net52),
    .X(_02156_));
 sky130_fd_sc_hd__a22o_1 _09953_ (.A1(_04268_),
    .A2(_01546_),
    .B1(_02156_),
    .B2(_01372_),
    .X(_02157_));
 sky130_fd_sc_hd__clkbuf_4 _09954_ (.A(_01546_),
    .X(_02158_));
 sky130_fd_sc_hd__nand4_2 _09955_ (.A(_04081_),
    .B(_01339_),
    .C(_02158_),
    .D(_02156_),
    .Y(_02159_));
 sky130_fd_sc_hd__and2_1 _09956_ (.A(_02157_),
    .B(_02159_),
    .X(_02161_));
 sky130_fd_sc_hd__xnor2_1 _09957_ (.A(_02155_),
    .B(_02161_),
    .Y(_02162_));
 sky130_fd_sc_hd__nor2_1 _09958_ (.A(_02154_),
    .B(_02162_),
    .Y(_02163_));
 sky130_fd_sc_hd__nand2_1 _09959_ (.A(_02154_),
    .B(_02162_),
    .Y(_02164_));
 sky130_fd_sc_hd__and2b_1 _09960_ (.A_N(_02163_),
    .B(_02164_),
    .X(_02165_));
 sky130_fd_sc_hd__a21o_1 _09961_ (.A1(_01661_),
    .A2(_01929_),
    .B1(_01928_),
    .X(_02166_));
 sky130_fd_sc_hd__xor2_2 _09962_ (.A(_02165_),
    .B(_02166_),
    .X(_02167_));
 sky130_fd_sc_hd__clkbuf_4 _09963_ (.A(net54),
    .X(_02168_));
 sky130_fd_sc_hd__clkbuf_4 _09964_ (.A(_02168_),
    .X(_02169_));
 sky130_fd_sc_hd__a22o_1 _09965_ (.A1(_02051_),
    .A2(_01934_),
    .B1(_02169_),
    .B2(_00453_),
    .X(_02170_));
 sky130_fd_sc_hd__and3_1 _09966_ (.A(_03576_),
    .B(_00989_),
    .C(net54),
    .X(_02172_));
 sky130_fd_sc_hd__nand2_1 _09967_ (.A(_01934_),
    .B(_02172_),
    .Y(_02173_));
 sky130_fd_sc_hd__nand2_1 _09968_ (.A(_02170_),
    .B(_02173_),
    .Y(_02174_));
 sky130_fd_sc_hd__xnor2_1 _09969_ (.A(_02167_),
    .B(_02174_),
    .Y(_02175_));
 sky130_fd_sc_hd__a22oi_1 _09970_ (.A1(_02171_),
    .A2(_01060_),
    .B1(_01413_),
    .B2(_02259_),
    .Y(_02176_));
 sky130_fd_sc_hd__and4_1 _09971_ (.A(_02105_),
    .B(_02149_),
    .C(_01058_),
    .D(_01411_),
    .X(_02177_));
 sky130_fd_sc_hd__nor2_1 _09972_ (.A(_02176_),
    .B(_02177_),
    .Y(_02178_));
 sky130_fd_sc_hd__xnor2_1 _09973_ (.A(_02175_),
    .B(_02178_),
    .Y(_02179_));
 sky130_fd_sc_hd__or2_2 _09974_ (.A(_02153_),
    .B(_02179_),
    .X(_02180_));
 sky130_fd_sc_hd__nand2_1 _09975_ (.A(_02153_),
    .B(_02179_),
    .Y(_02181_));
 sky130_fd_sc_hd__nand2_1 _09976_ (.A(_02180_),
    .B(_02181_),
    .Y(_02183_));
 sky130_fd_sc_hd__inv_2 _09977_ (.A(_02183_),
    .Y(_02184_));
 sky130_fd_sc_hd__or2b_1 _09978_ (.A(_01891_),
    .B_N(_01898_),
    .X(_02185_));
 sky130_fd_sc_hd__a31o_1 _09979_ (.A1(_06637_),
    .A2(_01400_),
    .A3(_01892_),
    .B1(_01893_),
    .X(_02186_));
 sky130_fd_sc_hd__clkbuf_4 _09980_ (.A(_01664_),
    .X(_02187_));
 sky130_fd_sc_hd__clkbuf_4 _09981_ (.A(_02187_),
    .X(_02188_));
 sky130_fd_sc_hd__clkbuf_4 _09982_ (.A(_01505_),
    .X(_02189_));
 sky130_fd_sc_hd__clkbuf_4 _09983_ (.A(_02189_),
    .X(_02190_));
 sky130_fd_sc_hd__a22oi_1 _09984_ (.A1(_06637_),
    .A2(_02188_),
    .B1(_02190_),
    .B2(_06937_),
    .Y(_02191_));
 sky130_fd_sc_hd__and4_1 _09985_ (.A(_06937_),
    .B(_06637_),
    .C(_02187_),
    .D(_02189_),
    .X(_02192_));
 sky130_fd_sc_hd__nor2_1 _09986_ (.A(_02191_),
    .B(_02192_),
    .Y(_02194_));
 sky130_fd_sc_hd__and2_1 _09987_ (.A(_02186_),
    .B(_02194_),
    .X(_02195_));
 sky130_fd_sc_hd__nor2_1 _09988_ (.A(_02186_),
    .B(_02194_),
    .Y(_02196_));
 sky130_fd_sc_hd__nor2_1 _09989_ (.A(_02195_),
    .B(_02196_),
    .Y(_02197_));
 sky130_fd_sc_hd__xnor2_1 _09990_ (.A(_02185_),
    .B(_02197_),
    .Y(_02198_));
 sky130_fd_sc_hd__a31o_1 _09991_ (.A1(_01535_),
    .A2(_01676_),
    .A3(_01902_),
    .B1(_01900_),
    .X(_02199_));
 sky130_fd_sc_hd__nor2_1 _09992_ (.A(_02198_),
    .B(_02199_),
    .Y(_02200_));
 sky130_fd_sc_hd__and2_1 _09993_ (.A(_02198_),
    .B(_02199_),
    .X(_02201_));
 sky130_fd_sc_hd__nor2_1 _09994_ (.A(_02200_),
    .B(_02201_),
    .Y(_02202_));
 sky130_fd_sc_hd__or2_1 _09995_ (.A(_01904_),
    .B(_02202_),
    .X(_02203_));
 sky130_fd_sc_hd__nand2_1 _09996_ (.A(_01904_),
    .B(_02202_),
    .Y(_02205_));
 sky130_fd_sc_hd__nand2_1 _09997_ (.A(_02203_),
    .B(_02205_),
    .Y(_02206_));
 sky130_fd_sc_hd__a21o_1 _09998_ (.A1(_01912_),
    .A2(_01915_),
    .B1(_01910_),
    .X(_02207_));
 sky130_fd_sc_hd__xnor2_2 _09999_ (.A(_02206_),
    .B(_02207_),
    .Y(_02208_));
 sky130_fd_sc_hd__xnor2_1 _10000_ (.A(_02184_),
    .B(_02208_),
    .Y(_02209_));
 sky130_fd_sc_hd__a21bo_1 _10001_ (.A1(_01869_),
    .A2(_01885_),
    .B1_N(_01887_),
    .X(_02210_));
 sky130_fd_sc_hd__nand2_1 _10002_ (.A(_01872_),
    .B(_01878_),
    .Y(_02211_));
 sky130_fd_sc_hd__a31o_1 _10003_ (.A1(_05181_),
    .A2(_04037_),
    .A3(_01876_),
    .B1(_01874_),
    .X(_02212_));
 sky130_fd_sc_hd__a22o_1 _10004_ (.A1(_04598_),
    .A2(_00612_),
    .B1(_00613_),
    .B2(_05192_),
    .X(_02213_));
 sky130_fd_sc_hd__nand4_1 _10005_ (.A(_05203_),
    .B(_04598_),
    .C(_00782_),
    .D(_00613_),
    .Y(_02214_));
 sky130_fd_sc_hd__and2_1 _10006_ (.A(_02213_),
    .B(_02214_),
    .X(_02216_));
 sky130_fd_sc_hd__xnor2_1 _10007_ (.A(_02212_),
    .B(_02216_),
    .Y(_02217_));
 sky130_fd_sc_hd__nor2_1 _10008_ (.A(_02211_),
    .B(_02217_),
    .Y(_02218_));
 sky130_fd_sc_hd__nand2_1 _10009_ (.A(_02211_),
    .B(_02217_),
    .Y(_02219_));
 sky130_fd_sc_hd__and2b_1 _10010_ (.A_N(_02218_),
    .B(_02219_),
    .X(_02220_));
 sky130_fd_sc_hd__a21o_1 _10011_ (.A1(_01709_),
    .A2(_01881_),
    .B1(_01880_),
    .X(_02221_));
 sky130_fd_sc_hd__xor2_2 _10012_ (.A(_02220_),
    .B(_02221_),
    .X(_02222_));
 sky130_fd_sc_hd__a22o_1 _10013_ (.A1(_03015_),
    .A2(_00458_),
    .B1(_00608_),
    .B2(_00388_),
    .X(_02223_));
 sky130_fd_sc_hd__and3_1 _10014_ (.A(_00366_),
    .B(_02971_),
    .C(net46),
    .X(_02224_));
 sky130_fd_sc_hd__nand2_1 _10015_ (.A(_00459_),
    .B(_02224_),
    .Y(_02225_));
 sky130_fd_sc_hd__nand2_1 _10016_ (.A(_02223_),
    .B(_02225_),
    .Y(_02227_));
 sky130_fd_sc_hd__xnor2_1 _10017_ (.A(_02222_),
    .B(_02227_),
    .Y(_02228_));
 sky130_fd_sc_hd__a22oi_1 _10018_ (.A1(_04939_),
    .A2(_00376_),
    .B1(_00379_),
    .B2(_04917_),
    .Y(_02229_));
 sky130_fd_sc_hd__and4_1 _10019_ (.A(_04862_),
    .B(_04873_),
    .C(_04037_),
    .D(_04059_),
    .X(_02230_));
 sky130_fd_sc_hd__nor2_1 _10020_ (.A(_02229_),
    .B(_02230_),
    .Y(_02231_));
 sky130_fd_sc_hd__xnor2_1 _10021_ (.A(_02228_),
    .B(_02231_),
    .Y(_02232_));
 sky130_fd_sc_hd__or2_4 _10022_ (.A(_02210_),
    .B(_02232_),
    .X(_02233_));
 sky130_fd_sc_hd__nand2_1 _10023_ (.A(_02210_),
    .B(_02232_),
    .Y(_02234_));
 sky130_fd_sc_hd__nand2_2 _10024_ (.A(_02233_),
    .B(_02234_),
    .Y(_02235_));
 sky130_fd_sc_hd__xnor2_2 _10025_ (.A(_02209_),
    .B(_02235_),
    .Y(_02236_));
 sky130_fd_sc_hd__a21o_1 _10026_ (.A1(_01916_),
    .A2(_01939_),
    .B1(_01889_),
    .X(_02238_));
 sky130_fd_sc_hd__o21a_1 _10027_ (.A1(_01916_),
    .A2(_01939_),
    .B1(_02238_),
    .X(_02239_));
 sky130_fd_sc_hd__xnor2_2 _10028_ (.A(_02236_),
    .B(_02239_),
    .Y(_02240_));
 sky130_fd_sc_hd__o31ai_4 _10029_ (.A1(_02152_),
    .A2(_01948_),
    .A3(_01949_),
    .B1(_02240_),
    .Y(_02241_));
 sky130_fd_sc_hd__o41a_2 _10030_ (.A1(_02152_),
    .A2(_01948_),
    .A3(_01949_),
    .A4(_02240_),
    .B1(_02241_),
    .X(_02242_));
 sky130_fd_sc_hd__inv_2 _10031_ (.A(_01753_),
    .Y(_02243_));
 sky130_fd_sc_hd__o211a_2 _10032_ (.A1(_01489_),
    .A2(_01488_),
    .B1(_02243_),
    .C1(_01867_),
    .X(_02244_));
 sky130_fd_sc_hd__o21ba_1 _10033_ (.A1(_01735_),
    .A2(_01851_),
    .B1_N(_01850_),
    .X(_02245_));
 sky130_fd_sc_hd__buf_4 _10034_ (.A(_00843_),
    .X(_02246_));
 sky130_fd_sc_hd__clkbuf_4 _10035_ (.A(_00859_),
    .X(_02247_));
 sky130_fd_sc_hd__clkbuf_4 _10036_ (.A(_00844_),
    .X(_02249_));
 sky130_fd_sc_hd__a22oi_1 _10037_ (.A1(_02246_),
    .A2(_01473_),
    .B1(_02247_),
    .B2(_02249_),
    .Y(_02250_));
 sky130_fd_sc_hd__and4_1 _10038_ (.A(_02246_),
    .B(_02249_),
    .C(_01473_),
    .D(_02247_),
    .X(_02251_));
 sky130_fd_sc_hd__nor2_1 _10039_ (.A(_02250_),
    .B(_02251_),
    .Y(_02252_));
 sky130_fd_sc_hd__o21a_1 _10040_ (.A1(_01841_),
    .A2(_01844_),
    .B1(_02252_),
    .X(_02253_));
 sky130_fd_sc_hd__nor3_1 _10041_ (.A(_01841_),
    .B(_01844_),
    .C(_02252_),
    .Y(_02254_));
 sky130_fd_sc_hd__nor2_1 _10042_ (.A(_02253_),
    .B(_02254_),
    .Y(_02255_));
 sky130_fd_sc_hd__and2_1 _10043_ (.A(_01847_),
    .B(_02255_),
    .X(_02256_));
 sky130_fd_sc_hd__nor2_1 _10044_ (.A(_01847_),
    .B(_02255_),
    .Y(_02257_));
 sky130_fd_sc_hd__nor2_1 _10045_ (.A(_02256_),
    .B(_02257_),
    .Y(_02258_));
 sky130_fd_sc_hd__and2b_1 _10046_ (.A_N(_02245_),
    .B(_02258_),
    .X(_02260_));
 sky130_fd_sc_hd__and2b_1 _10047_ (.A_N(_02258_),
    .B(_02245_),
    .X(_02261_));
 sky130_fd_sc_hd__nor2_1 _10048_ (.A(_02260_),
    .B(_02261_),
    .Y(_02262_));
 sky130_fd_sc_hd__nand2_1 _10049_ (.A(_01855_),
    .B(_02262_),
    .Y(_02263_));
 sky130_fd_sc_hd__or2_1 _10050_ (.A(_01855_),
    .B(_02262_),
    .X(_02264_));
 sky130_fd_sc_hd__nand2_1 _10051_ (.A(_02263_),
    .B(_02264_),
    .Y(_02265_));
 sky130_fd_sc_hd__o21bai_2 _10052_ (.A1(_01859_),
    .A2(_01865_),
    .B1_N(_02265_),
    .Y(_02266_));
 sky130_fd_sc_hd__or3b_1 _10053_ (.A(_01859_),
    .B(_01865_),
    .C_N(_02265_),
    .X(_02267_));
 sky130_fd_sc_hd__nand2_2 _10054_ (.A(_02266_),
    .B(_02267_),
    .Y(_02268_));
 sky130_fd_sc_hd__xnor2_4 _10055_ (.A(_02244_),
    .B(_02268_),
    .Y(_02269_));
 sky130_fd_sc_hd__xor2_2 _10056_ (.A(_02242_),
    .B(_02269_),
    .X(_02271_));
 sky130_fd_sc_hd__xnor2_4 _10057_ (.A(_02151_),
    .B(_02271_),
    .Y(_02272_));
 sky130_fd_sc_hd__xor2_4 _10058_ (.A(_02055_),
    .B(_02272_),
    .X(_02273_));
 sky130_fd_sc_hd__xor2_4 _10059_ (.A(_02052_),
    .B(_02273_),
    .X(_02274_));
 sky130_fd_sc_hd__and2_1 _10060_ (.A(_01837_),
    .B(_02045_),
    .X(_02275_));
 sky130_fd_sc_hd__a21oi_1 _10061_ (.A1(_01833_),
    .A2(_01835_),
    .B1(_02044_),
    .Y(_02276_));
 sky130_fd_sc_hd__a41o_1 _10062_ (.A1(_01646_),
    .A2(_01643_),
    .A3(_01837_),
    .A4(_02045_),
    .B1(_02276_),
    .X(_02277_));
 sky130_fd_sc_hd__a41o_2 _10063_ (.A1(_01433_),
    .A2(_01437_),
    .A3(_01636_),
    .A4(_02275_),
    .B1(_02277_),
    .X(_02278_));
 sky130_fd_sc_hd__xor2_2 _10064_ (.A(_02274_),
    .B(_02278_),
    .X(net86));
 sky130_fd_sc_hd__nor2_2 _10065_ (.A(_02055_),
    .B(_02272_),
    .Y(_02279_));
 sky130_fd_sc_hd__nand2_1 _10066_ (.A(_01752_),
    .B(_01867_),
    .Y(_02281_));
 sky130_fd_sc_hd__nor2_1 _10067_ (.A(_02268_),
    .B(_02281_),
    .Y(_02282_));
 sky130_fd_sc_hd__and3_1 _10068_ (.A(_02246_),
    .B(_02247_),
    .C(_01839_),
    .X(_02283_));
 sky130_fd_sc_hd__and2_1 _10069_ (.A(_02253_),
    .B(_02283_),
    .X(_02284_));
 sky130_fd_sc_hd__nor2_1 _10070_ (.A(_02253_),
    .B(_02283_),
    .Y(_02285_));
 sky130_fd_sc_hd__nor2_1 _10071_ (.A(_02284_),
    .B(_02285_),
    .Y(_02286_));
 sky130_fd_sc_hd__or3_1 _10072_ (.A(_02256_),
    .B(_02260_),
    .C(_02286_),
    .X(_02287_));
 sky130_fd_sc_hd__o21ai_1 _10073_ (.A1(_02256_),
    .A2(_02260_),
    .B1(_02286_),
    .Y(_02288_));
 sky130_fd_sc_hd__nand2_1 _10074_ (.A(_02287_),
    .B(_02288_),
    .Y(_02289_));
 sky130_fd_sc_hd__and3_1 _10075_ (.A(_02263_),
    .B(_02266_),
    .C(_02289_),
    .X(_02290_));
 sky130_fd_sc_hd__a21o_1 _10076_ (.A1(_02263_),
    .A2(_02266_),
    .B1(_02289_),
    .X(_02292_));
 sky130_fd_sc_hd__and2b_1 _10077_ (.A_N(_02290_),
    .B(_02292_),
    .X(_02293_));
 sky130_fd_sc_hd__and2_1 _10078_ (.A(_02282_),
    .B(_02293_),
    .X(_02294_));
 sky130_fd_sc_hd__nor2_1 _10079_ (.A(_02282_),
    .B(_02293_),
    .Y(_02295_));
 sky130_fd_sc_hd__a2111o_1 _10080_ (.A1(_01443_),
    .A2(_01444_),
    .B1(_02294_),
    .C1(_02295_),
    .D1(_01486_),
    .X(_02296_));
 sky130_fd_sc_hd__inv_2 _10081_ (.A(_02293_),
    .Y(_02297_));
 sky130_fd_sc_hd__a311o_1 _10082_ (.A1(_00991_),
    .A2(_01356_),
    .A3(_01756_),
    .B1(_01757_),
    .C1(_02297_),
    .X(_02298_));
 sky130_fd_sc_hd__or2b_1 _10083_ (.A(_02236_),
    .B_N(_02239_),
    .X(_02299_));
 sky130_fd_sc_hd__or2b_1 _10084_ (.A(_02167_),
    .B_N(_02174_),
    .X(_02300_));
 sky130_fd_sc_hd__a32o_1 _10085_ (.A1(_02167_),
    .A2(_02170_),
    .A3(_02173_),
    .B1(_02300_),
    .B2(_02178_),
    .X(_02301_));
 sky130_fd_sc_hd__and2_1 _10086_ (.A(_02155_),
    .B(_02161_),
    .X(_02303_));
 sky130_fd_sc_hd__buf_2 _10087_ (.A(_02156_),
    .X(_02304_));
 sky130_fd_sc_hd__clkbuf_4 _10088_ (.A(_02304_),
    .X(_02305_));
 sky130_fd_sc_hd__clkbuf_4 _10089_ (.A(_02158_),
    .X(_02306_));
 sky130_fd_sc_hd__nand2_1 _10090_ (.A(_01383_),
    .B(_02306_),
    .Y(_02307_));
 sky130_fd_sc_hd__and3_2 _10091_ (.A(_01350_),
    .B(_02305_),
    .C(_02307_),
    .X(_02308_));
 sky130_fd_sc_hd__xor2_2 _10092_ (.A(_02303_),
    .B(_02308_),
    .X(_02309_));
 sky130_fd_sc_hd__a21o_1 _10093_ (.A1(_02165_),
    .A2(_02166_),
    .B1(_02163_),
    .X(_02310_));
 sky130_fd_sc_hd__xnor2_2 _10094_ (.A(_02309_),
    .B(_02310_),
    .Y(_02311_));
 sky130_fd_sc_hd__buf_2 _10095_ (.A(net56),
    .X(_02312_));
 sky130_fd_sc_hd__a22o_1 _10096_ (.A1(_00989_),
    .A2(net54),
    .B1(_02312_),
    .B2(_03576_),
    .X(_02314_));
 sky130_fd_sc_hd__a21bo_1 _10097_ (.A1(_02312_),
    .A2(_02172_),
    .B1_N(_02314_),
    .X(_02315_));
 sky130_fd_sc_hd__nand2_1 _10098_ (.A(_04081_),
    .B(net53),
    .Y(_02316_));
 sky130_fd_sc_hd__xor2_1 _10099_ (.A(_02315_),
    .B(_02316_),
    .X(_02317_));
 sky130_fd_sc_hd__and3_1 _10100_ (.A(_01933_),
    .B(_02172_),
    .C(_02317_),
    .X(_02318_));
 sky130_fd_sc_hd__a21oi_1 _10101_ (.A1(_01934_),
    .A2(_02172_),
    .B1(_02317_),
    .Y(_02319_));
 sky130_fd_sc_hd__or2_1 _10102_ (.A(_02318_),
    .B(_02319_),
    .X(_02320_));
 sky130_fd_sc_hd__xnor2_1 _10103_ (.A(_02311_),
    .B(_02320_),
    .Y(_02321_));
 sky130_fd_sc_hd__a22oi_1 _10104_ (.A1(_00650_),
    .A2(_01410_),
    .B1(_02158_),
    .B2(_02105_),
    .Y(_02322_));
 sky130_fd_sc_hd__and4_1 _10105_ (.A(_00628_),
    .B(_05742_),
    .C(net50),
    .D(_01545_),
    .X(_02323_));
 sky130_fd_sc_hd__o2bb2a_1 _10106_ (.A1_N(_05588_),
    .A2_N(_01058_),
    .B1(_02322_),
    .B2(_02323_),
    .X(_02325_));
 sky130_fd_sc_hd__a22o_1 _10107_ (.A1(_05742_),
    .A2(net50),
    .B1(_01546_),
    .B2(_00628_),
    .X(_02326_));
 sky130_fd_sc_hd__and4b_1 _10108_ (.A_N(_02323_),
    .B(_01058_),
    .C(_05577_),
    .D(_02326_),
    .X(_02327_));
 sky130_fd_sc_hd__nor2_1 _10109_ (.A(_02325_),
    .B(_02327_),
    .Y(_02328_));
 sky130_fd_sc_hd__and2_1 _10110_ (.A(_02177_),
    .B(_02328_),
    .X(_02329_));
 sky130_fd_sc_hd__nor2_1 _10111_ (.A(_02177_),
    .B(_02328_),
    .Y(_02330_));
 sky130_fd_sc_hd__nor2_1 _10112_ (.A(_02329_),
    .B(_02330_),
    .Y(_02331_));
 sky130_fd_sc_hd__xnor2_2 _10113_ (.A(_02321_),
    .B(_02331_),
    .Y(_02332_));
 sky130_fd_sc_hd__xnor2_2 _10114_ (.A(_02301_),
    .B(_02332_),
    .Y(_02333_));
 sky130_fd_sc_hd__xor2_2 _10115_ (.A(_02180_),
    .B(_02333_),
    .X(_02334_));
 sky130_fd_sc_hd__and2b_1 _10116_ (.A_N(_02185_),
    .B(_02197_),
    .X(_02336_));
 sky130_fd_sc_hd__nand2_1 _10117_ (.A(_06937_),
    .B(_02188_),
    .Y(_02337_));
 sky130_fd_sc_hd__and3_1 _10118_ (.A(_06637_),
    .B(_02190_),
    .C(_02337_),
    .X(_02338_));
 sky130_fd_sc_hd__xor2_1 _10119_ (.A(_02195_),
    .B(_02338_),
    .X(_02339_));
 sky130_fd_sc_hd__nor3_1 _10120_ (.A(_02336_),
    .B(_02201_),
    .C(_02339_),
    .Y(_02340_));
 sky130_fd_sc_hd__o21a_1 _10121_ (.A1(_02336_),
    .A2(_02201_),
    .B1(_02339_),
    .X(_02341_));
 sky130_fd_sc_hd__nor2_2 _10122_ (.A(_02340_),
    .B(_02341_),
    .Y(_02342_));
 sky130_fd_sc_hd__o21a_1 _10123_ (.A1(_01904_),
    .A2(_01910_),
    .B1(_02202_),
    .X(_02343_));
 sky130_fd_sc_hd__a31oi_4 _10124_ (.A1(_01912_),
    .A2(_01915_),
    .A3(_02203_),
    .B1(_02343_),
    .Y(_02344_));
 sky130_fd_sc_hd__xnor2_2 _10125_ (.A(_02342_),
    .B(_02344_),
    .Y(_02345_));
 sky130_fd_sc_hd__xnor2_1 _10126_ (.A(_02334_),
    .B(_02345_),
    .Y(_02347_));
 sky130_fd_sc_hd__or2b_1 _10127_ (.A(_02222_),
    .B_N(_02227_),
    .X(_02348_));
 sky130_fd_sc_hd__a32o_2 _10128_ (.A1(_02222_),
    .A2(_02223_),
    .A3(_02225_),
    .B1(_02348_),
    .B2(_02231_),
    .X(_02349_));
 sky130_fd_sc_hd__and2_1 _10129_ (.A(_02212_),
    .B(_02216_),
    .X(_02350_));
 sky130_fd_sc_hd__nand2_1 _10130_ (.A(_00094_),
    .B(_00784_),
    .Y(_02351_));
 sky130_fd_sc_hd__and3_1 _10131_ (.A(_00151_),
    .B(_01517_),
    .C(_02351_),
    .X(_02352_));
 sky130_fd_sc_hd__xor2_2 _10132_ (.A(_02350_),
    .B(_02352_),
    .X(_02353_));
 sky130_fd_sc_hd__a21o_1 _10133_ (.A1(_02220_),
    .A2(_02221_),
    .B1(_02218_),
    .X(_02354_));
 sky130_fd_sc_hd__xnor2_2 _10134_ (.A(_02353_),
    .B(_02354_),
    .Y(_02355_));
 sky130_fd_sc_hd__a22o_1 _10135_ (.A1(_02971_),
    .A2(net46),
    .B1(_01368_),
    .B2(_00366_),
    .X(_02356_));
 sky130_fd_sc_hd__a21bo_1 _10136_ (.A1(_01506_),
    .A2(_02224_),
    .B1_N(_02356_),
    .X(_02358_));
 sky130_fd_sc_hd__nand2_1 _10137_ (.A(_05203_),
    .B(net45),
    .Y(_02359_));
 sky130_fd_sc_hd__xor2_1 _10138_ (.A(_02358_),
    .B(_02359_),
    .X(_02360_));
 sky130_fd_sc_hd__and3_1 _10139_ (.A(_00457_),
    .B(_02224_),
    .C(_02360_),
    .X(_02361_));
 sky130_fd_sc_hd__a21oi_1 _10140_ (.A1(_00458_),
    .A2(_02224_),
    .B1(_02360_),
    .Y(_02362_));
 sky130_fd_sc_hd__or2_2 _10141_ (.A(_02361_),
    .B(_02362_),
    .X(_02363_));
 sky130_fd_sc_hd__xnor2_2 _10142_ (.A(_02355_),
    .B(_02363_),
    .Y(_02364_));
 sky130_fd_sc_hd__a22oi_1 _10143_ (.A1(_04862_),
    .A2(_00373_),
    .B1(_00782_),
    .B2(_04873_),
    .Y(_02365_));
 sky130_fd_sc_hd__and4_1 _10144_ (.A(_04851_),
    .B(net4),
    .C(_04015_),
    .D(_00780_),
    .X(_02366_));
 sky130_fd_sc_hd__o2bb2a_1 _10145_ (.A1_N(_05027_),
    .A2_N(_04048_),
    .B1(_02365_),
    .B2(_02366_),
    .X(_02367_));
 sky130_fd_sc_hd__a22o_1 _10146_ (.A1(_04851_),
    .A2(_04015_),
    .B1(_00780_),
    .B2(net4),
    .X(_02369_));
 sky130_fd_sc_hd__and4b_1 _10147_ (.A_N(_02366_),
    .B(_04048_),
    .C(_05027_),
    .D(_02369_),
    .X(_02370_));
 sky130_fd_sc_hd__nor2_1 _10148_ (.A(_02367_),
    .B(_02370_),
    .Y(_02371_));
 sky130_fd_sc_hd__and2_1 _10149_ (.A(_02230_),
    .B(_02371_),
    .X(_02372_));
 sky130_fd_sc_hd__nor2_1 _10150_ (.A(_02230_),
    .B(_02371_),
    .Y(_02373_));
 sky130_fd_sc_hd__nor2_2 _10151_ (.A(_02372_),
    .B(_02373_),
    .Y(_02374_));
 sky130_fd_sc_hd__xnor2_4 _10152_ (.A(_02364_),
    .B(_02374_),
    .Y(_02375_));
 sky130_fd_sc_hd__xnor2_4 _10153_ (.A(_02349_),
    .B(_02375_),
    .Y(_02376_));
 sky130_fd_sc_hd__xnor2_4 _10154_ (.A(_02233_),
    .B(_02376_),
    .Y(_02377_));
 sky130_fd_sc_hd__xnor2_1 _10155_ (.A(_02347_),
    .B(_02377_),
    .Y(_02378_));
 sky130_fd_sc_hd__a21bo_1 _10156_ (.A1(_02184_),
    .A2(_02208_),
    .B1_N(_02235_),
    .X(_02380_));
 sky130_fd_sc_hd__o21ai_1 _10157_ (.A1(_02184_),
    .A2(_02208_),
    .B1(_02380_),
    .Y(_02381_));
 sky130_fd_sc_hd__or2_2 _10158_ (.A(_02378_),
    .B(_02381_),
    .X(_02382_));
 sky130_fd_sc_hd__nand2_1 _10159_ (.A(_02378_),
    .B(_02381_),
    .Y(_02383_));
 sky130_fd_sc_hd__nand2_1 _10160_ (.A(_02382_),
    .B(_02383_),
    .Y(_02384_));
 sky130_fd_sc_hd__a21o_1 _10161_ (.A1(_02299_),
    .A2(_02241_),
    .B1(_02384_),
    .X(_02385_));
 sky130_fd_sc_hd__nand3_1 _10162_ (.A(_02299_),
    .B(_02241_),
    .C(_02384_),
    .Y(_02386_));
 sky130_fd_sc_hd__nand2_1 _10163_ (.A(_02385_),
    .B(_02386_),
    .Y(_02387_));
 sky130_fd_sc_hd__a21o_1 _10164_ (.A1(_02296_),
    .A2(_02298_),
    .B1(_02387_),
    .X(_02388_));
 sky130_fd_sc_hd__nand3_2 _10165_ (.A(_02387_),
    .B(_02296_),
    .C(_02298_),
    .Y(_02389_));
 sky130_fd_sc_hd__or2b_1 _10166_ (.A(_02145_),
    .B_N(_02147_),
    .X(_02391_));
 sky130_fd_sc_hd__a21bo_1 _10167_ (.A1(_02074_),
    .A2(_02080_),
    .B1_N(_02075_),
    .X(_02392_));
 sky130_fd_sc_hd__and3_1 _10168_ (.A(_02063_),
    .B(_02064_),
    .C(_02065_),
    .X(_02393_));
 sky130_fd_sc_hd__and3_1 _10169_ (.A(_06965_),
    .B(_00741_),
    .C(_02014_),
    .X(_02394_));
 sky130_fd_sc_hd__and2_1 _10170_ (.A(_02393_),
    .B(_02394_),
    .X(_02395_));
 sky130_fd_sc_hd__nor2_1 _10171_ (.A(_02393_),
    .B(_02394_),
    .Y(_02396_));
 sky130_fd_sc_hd__nor2_1 _10172_ (.A(_02395_),
    .B(_02396_),
    .Y(_02397_));
 sky130_fd_sc_hd__a21o_1 _10173_ (.A1(_02069_),
    .A2(_02071_),
    .B1(_02068_),
    .X(_02398_));
 sky130_fd_sc_hd__xnor2_2 _10174_ (.A(_02397_),
    .B(_02398_),
    .Y(_02399_));
 sky130_fd_sc_hd__a22o_1 _10175_ (.A1(_00101_),
    .A2(_03685_),
    .B1(_03718_),
    .B2(net37),
    .X(_02400_));
 sky130_fd_sc_hd__inv_2 _10176_ (.A(_02400_),
    .Y(_02402_));
 sky130_fd_sc_hd__and4_1 _10177_ (.A(_00101_),
    .B(_06733_),
    .C(_03685_),
    .D(_00423_),
    .X(_02403_));
 sky130_fd_sc_hd__o2bb2a_1 _10178_ (.A1_N(_06744_),
    .A2_N(_03773_),
    .B1(_02402_),
    .B2(_02403_),
    .X(_02404_));
 sky130_fd_sc_hd__and4b_1 _10179_ (.A_N(_02403_),
    .B(_03894_),
    .C(_06744_),
    .D(_02400_),
    .X(_02405_));
 sky130_fd_sc_hd__or2_1 _10180_ (.A(_02404_),
    .B(_02405_),
    .X(_02406_));
 sky130_fd_sc_hd__or2_2 _10181_ (.A(_02060_),
    .B(_02406_),
    .X(_02407_));
 sky130_fd_sc_hd__nand2_1 _10182_ (.A(_02060_),
    .B(_02406_),
    .Y(_02408_));
 sky130_fd_sc_hd__nand2_2 _10183_ (.A(_02407_),
    .B(_02408_),
    .Y(_02409_));
 sky130_fd_sc_hd__xor2_2 _10184_ (.A(_02399_),
    .B(_02409_),
    .X(_02410_));
 sky130_fd_sc_hd__a22o_1 _10185_ (.A1(_06821_),
    .A2(net13),
    .B1(_00730_),
    .B2(_03499_),
    .X(_02411_));
 sky130_fd_sc_hd__inv_2 _10186_ (.A(_02411_),
    .Y(_02413_));
 sky130_fd_sc_hd__and4_1 _10187_ (.A(_03499_),
    .B(_06821_),
    .C(net13),
    .D(_00730_),
    .X(_02414_));
 sky130_fd_sc_hd__o2bb2a_1 _10188_ (.A1_N(_00486_),
    .A2_N(_00734_),
    .B1(_02413_),
    .B2(_02414_),
    .X(_02415_));
 sky130_fd_sc_hd__and4b_1 _10189_ (.A_N(_02414_),
    .B(_00734_),
    .C(_00486_),
    .D(_02411_),
    .X(_02416_));
 sky130_fd_sc_hd__or2_1 _10190_ (.A(_02415_),
    .B(_02416_),
    .X(_02417_));
 sky130_fd_sc_hd__or2_1 _10191_ (.A(_02079_),
    .B(_02417_),
    .X(_02418_));
 sky130_fd_sc_hd__nand2_1 _10192_ (.A(_02079_),
    .B(_02417_),
    .Y(_02419_));
 sky130_fd_sc_hd__nand2_1 _10193_ (.A(_02418_),
    .B(_02419_),
    .Y(_02420_));
 sky130_fd_sc_hd__xnor2_2 _10194_ (.A(_02410_),
    .B(_02420_),
    .Y(_02421_));
 sky130_fd_sc_hd__xor2_2 _10195_ (.A(_02392_),
    .B(_02421_),
    .X(_02422_));
 sky130_fd_sc_hd__xor2_2 _10196_ (.A(_02082_),
    .B(_02422_),
    .X(_02424_));
 sky130_fd_sc_hd__and2b_1 _10197_ (.A_N(_02087_),
    .B(_02097_),
    .X(_02425_));
 sky130_fd_sc_hd__clkbuf_4 _10198_ (.A(_02088_),
    .X(_02426_));
 sky130_fd_sc_hd__clkbuf_4 _10199_ (.A(_02090_),
    .X(_02427_));
 sky130_fd_sc_hd__nand2_1 _10200_ (.A(_06450_),
    .B(_02427_),
    .Y(_02428_));
 sky130_fd_sc_hd__and3_1 _10201_ (.A(_06626_),
    .B(_02426_),
    .C(_02428_),
    .X(_02429_));
 sky130_fd_sc_hd__xor2_1 _10202_ (.A(_02095_),
    .B(_02429_),
    .X(_02430_));
 sky130_fd_sc_hd__nor3_1 _10203_ (.A(_02425_),
    .B(_02101_),
    .C(_02430_),
    .Y(_02431_));
 sky130_fd_sc_hd__o21a_1 _10204_ (.A1(_02425_),
    .A2(_02101_),
    .B1(_02430_),
    .X(_02432_));
 sky130_fd_sc_hd__nor2_1 _10205_ (.A(_02431_),
    .B(_02432_),
    .Y(_02433_));
 sky130_fd_sc_hd__o21a_1 _10206_ (.A1(_01995_),
    .A2(_02001_),
    .B1(_02102_),
    .X(_02435_));
 sky130_fd_sc_hd__a31oi_4 _10207_ (.A1(_02003_),
    .A2(_02005_),
    .A3(_02103_),
    .B1(_02435_),
    .Y(_02436_));
 sky130_fd_sc_hd__xnor2_2 _10208_ (.A(_02433_),
    .B(_02436_),
    .Y(_02437_));
 sky130_fd_sc_hd__xnor2_1 _10209_ (.A(_02424_),
    .B(_02437_),
    .Y(_02438_));
 sky130_fd_sc_hd__a21bo_1 _10210_ (.A1(_02130_),
    .A2(_02140_),
    .B1_N(_02131_),
    .X(_02439_));
 sky130_fd_sc_hd__and3_1 _10211_ (.A(_02115_),
    .B(_02118_),
    .C(_02121_),
    .X(_02440_));
 sky130_fd_sc_hd__and3_1 _10212_ (.A(_00157_),
    .B(_02120_),
    .C(_01966_),
    .X(_02441_));
 sky130_fd_sc_hd__and2_1 _10213_ (.A(_02440_),
    .B(_02441_),
    .X(_02442_));
 sky130_fd_sc_hd__nor2_1 _10214_ (.A(_02440_),
    .B(_02441_),
    .Y(_02443_));
 sky130_fd_sc_hd__nor2_1 _10215_ (.A(_02442_),
    .B(_02443_),
    .Y(_02444_));
 sky130_fd_sc_hd__a21o_1 _10216_ (.A1(_02125_),
    .A2(_02128_),
    .B1(_02124_),
    .X(_02446_));
 sky130_fd_sc_hd__xnor2_2 _10217_ (.A(_02444_),
    .B(_02446_),
    .Y(_02447_));
 sky130_fd_sc_hd__a22o_1 _10218_ (.A1(_05731_),
    .A2(_01177_),
    .B1(_01246_),
    .B2(_01000_),
    .X(_02448_));
 sky130_fd_sc_hd__inv_2 _10219_ (.A(_02448_),
    .Y(_02449_));
 sky130_fd_sc_hd__and4_1 _10220_ (.A(_05467_),
    .B(_01000_),
    .C(_01177_),
    .D(_01246_),
    .X(_02450_));
 sky130_fd_sc_hd__o2bb2a_1 _10221_ (.A1_N(_02029_),
    .A2_N(_01564_),
    .B1(_02449_),
    .B2(_02450_),
    .X(_02451_));
 sky130_fd_sc_hd__and4b_1 _10222_ (.A_N(_02450_),
    .B(_01564_),
    .C(_02029_),
    .D(_02448_),
    .X(_02452_));
 sky130_fd_sc_hd__or2_1 _10223_ (.A(_02451_),
    .B(_02452_),
    .X(_02453_));
 sky130_fd_sc_hd__or2_1 _10224_ (.A(_02113_),
    .B(_02453_),
    .X(_02454_));
 sky130_fd_sc_hd__nand2_1 _10225_ (.A(_02113_),
    .B(_02453_),
    .Y(_02455_));
 sky130_fd_sc_hd__nand2_1 _10226_ (.A(_02454_),
    .B(_02455_),
    .Y(_02457_));
 sky130_fd_sc_hd__xor2_1 _10227_ (.A(_02447_),
    .B(_02457_),
    .X(_02458_));
 sky130_fd_sc_hd__clkbuf_4 _10228_ (.A(net24),
    .X(_02459_));
 sky130_fd_sc_hd__a22o_1 _10229_ (.A1(_01394_),
    .A2(net21),
    .B1(net22),
    .B2(_01470_),
    .X(_02460_));
 sky130_fd_sc_hd__inv_2 _10230_ (.A(_02460_),
    .Y(_02461_));
 sky130_fd_sc_hd__and4_1 _10231_ (.A(_01306_),
    .B(_00672_),
    .C(net21),
    .D(net22),
    .X(_02462_));
 sky130_fd_sc_hd__o2bb2a_1 _10232_ (.A1_N(_00322_),
    .A2_N(_02459_),
    .B1(_02461_),
    .B2(_02462_),
    .X(_02463_));
 sky130_fd_sc_hd__and4b_1 _10233_ (.A_N(_02462_),
    .B(net24),
    .C(_00322_),
    .D(_02460_),
    .X(_02464_));
 sky130_fd_sc_hd__or2_1 _10234_ (.A(_02463_),
    .B(_02464_),
    .X(_02465_));
 sky130_fd_sc_hd__or2_1 _10235_ (.A(_02139_),
    .B(_02465_),
    .X(_02466_));
 sky130_fd_sc_hd__nand2_1 _10236_ (.A(_02139_),
    .B(_02465_),
    .Y(_02468_));
 sky130_fd_sc_hd__nand2_1 _10237_ (.A(_02466_),
    .B(_02468_),
    .Y(_02469_));
 sky130_fd_sc_hd__xnor2_2 _10238_ (.A(_02458_),
    .B(_02469_),
    .Y(_02470_));
 sky130_fd_sc_hd__xor2_2 _10239_ (.A(_02439_),
    .B(_02470_),
    .X(_02471_));
 sky130_fd_sc_hd__xnor2_2 _10240_ (.A(_02142_),
    .B(_02471_),
    .Y(_02472_));
 sky130_fd_sc_hd__xnor2_1 _10241_ (.A(_02438_),
    .B(_02472_),
    .Y(_02473_));
 sky130_fd_sc_hd__a21bo_1 _10242_ (.A1(_02086_),
    .A2(_02108_),
    .B1_N(_02144_),
    .X(_02474_));
 sky130_fd_sc_hd__o21ai_2 _10243_ (.A1(_02086_),
    .A2(_02108_),
    .B1(_02474_),
    .Y(_02475_));
 sky130_fd_sc_hd__nor2_1 _10244_ (.A(_02473_),
    .B(_02475_),
    .Y(_02476_));
 sky130_fd_sc_hd__and2_1 _10245_ (.A(_02473_),
    .B(_02475_),
    .X(_02477_));
 sky130_fd_sc_hd__or2_1 _10246_ (.A(_02476_),
    .B(_02477_),
    .X(_02479_));
 sky130_fd_sc_hd__a21oi_2 _10247_ (.A1(_02391_),
    .A2(_02150_),
    .B1(_02479_),
    .Y(_02480_));
 sky130_fd_sc_hd__and3_1 _10248_ (.A(_02391_),
    .B(_02150_),
    .C(_02479_),
    .X(_02481_));
 sky130_fd_sc_hd__or2_4 _10249_ (.A(_02480_),
    .B(_02481_),
    .X(_02482_));
 sky130_fd_sc_hd__a21o_1 _10250_ (.A1(_02388_),
    .A2(_02389_),
    .B1(_02482_),
    .X(_02483_));
 sky130_fd_sc_hd__nand3_2 _10251_ (.A(_02388_),
    .B(_02389_),
    .C(_02482_),
    .Y(_02484_));
 sky130_fd_sc_hd__nor2_1 _10252_ (.A(_02242_),
    .B(_02269_),
    .Y(_02485_));
 sky130_fd_sc_hd__a21oi_2 _10253_ (.A1(_02242_),
    .A2(_02269_),
    .B1(_02151_),
    .Y(_02486_));
 sky130_fd_sc_hd__a211oi_2 _10254_ (.A1(_02483_),
    .A2(_02484_),
    .B1(_02485_),
    .C1(_02486_),
    .Y(_02487_));
 sky130_fd_sc_hd__o211a_1 _10255_ (.A1(_02485_),
    .A2(_02486_),
    .B1(_02483_),
    .C1(_02484_),
    .X(_02488_));
 sky130_fd_sc_hd__or2_2 _10256_ (.A(_02487_),
    .B(_02488_),
    .X(_02490_));
 sky130_fd_sc_hd__xnor2_4 _10257_ (.A(_02279_),
    .B(_02490_),
    .Y(_02491_));
 sky130_fd_sc_hd__and2_2 _10258_ (.A(_02045_),
    .B(_02274_),
    .X(_02492_));
 sky130_fd_sc_hd__o21bai_1 _10259_ (.A1(_01833_),
    .A2(_02044_),
    .B1_N(_02052_),
    .Y(_02493_));
 sky130_fd_sc_hd__a32o_1 _10260_ (.A1(_02045_),
    .A2(_02049_),
    .A3(_02274_),
    .B1(_02493_),
    .B2(_02273_),
    .X(_02494_));
 sky130_fd_sc_hd__a31o_1 _10261_ (.A1(_01640_),
    .A2(_02046_),
    .A3(_02492_),
    .B1(_02494_),
    .X(_02495_));
 sky130_fd_sc_hd__xor2_1 _10262_ (.A(_02491_),
    .B(_02495_),
    .X(net88));
 sky130_fd_sc_hd__and4bb_2 _10263_ (.A_N(_02251_),
    .B_N(_02284_),
    .C(_02288_),
    .D(_02292_),
    .X(_02496_));
 sky130_fd_sc_hd__and2_1 _10264_ (.A(_01757_),
    .B(_02294_),
    .X(_02497_));
 sky130_fd_sc_hd__a41oi_4 _10265_ (.A1(_00991_),
    .A2(_01356_),
    .A3(_01756_),
    .A4(_02294_),
    .B1(_02497_),
    .Y(_02498_));
 sky130_fd_sc_hd__inv_2 _10266_ (.A(_02342_),
    .Y(_02500_));
 sky130_fd_sc_hd__a211oi_2 _10267_ (.A1(_02195_),
    .A2(_02338_),
    .B1(_02341_),
    .C1(_02192_),
    .Y(_02501_));
 sky130_fd_sc_hd__o21ai_4 _10268_ (.A1(_02500_),
    .A2(_02344_),
    .B1(_02501_),
    .Y(_02502_));
 sky130_fd_sc_hd__o21ba_1 _10269_ (.A1(_02311_),
    .A2(_02320_),
    .B1_N(_02331_),
    .X(_02503_));
 sky130_fd_sc_hd__a21o_1 _10270_ (.A1(_02311_),
    .A2(_02320_),
    .B1(_02503_),
    .X(_02504_));
 sky130_fd_sc_hd__nand2_1 _10271_ (.A(_02303_),
    .B(_02308_),
    .Y(_02505_));
 sky130_fd_sc_hd__nand2_1 _10272_ (.A(_02309_),
    .B(_02310_),
    .Y(_02506_));
 sky130_fd_sc_hd__and3_1 _10273_ (.A(_03576_),
    .B(_00989_),
    .C(_02312_),
    .X(_02507_));
 sky130_fd_sc_hd__a22o_1 _10274_ (.A1(_00989_),
    .A2(_02312_),
    .B1(net57),
    .B2(_03576_),
    .X(_02508_));
 sky130_fd_sc_hd__a21bo_1 _10275_ (.A1(net57),
    .A2(_02507_),
    .B1_N(_02508_),
    .X(_02509_));
 sky130_fd_sc_hd__nand2_1 _10276_ (.A(_04081_),
    .B(net54),
    .Y(_02511_));
 sky130_fd_sc_hd__xor2_1 _10277_ (.A(_02509_),
    .B(_02511_),
    .X(_02512_));
 sky130_fd_sc_hd__a32o_1 _10278_ (.A1(_01372_),
    .A2(net53),
    .A3(_02314_),
    .B1(_02172_),
    .B2(_02312_),
    .X(_02513_));
 sky130_fd_sc_hd__nand2_1 _10279_ (.A(_01339_),
    .B(net53),
    .Y(_02514_));
 sky130_fd_sc_hd__xnor2_1 _10280_ (.A(_02513_),
    .B(_02514_),
    .Y(_02515_));
 sky130_fd_sc_hd__xor2_1 _10281_ (.A(_02512_),
    .B(_02515_),
    .X(_02516_));
 sky130_fd_sc_hd__nand2_1 _10282_ (.A(_02318_),
    .B(_02516_),
    .Y(_02517_));
 sky130_fd_sc_hd__or2_1 _10283_ (.A(_02318_),
    .B(_02516_),
    .X(_02518_));
 sky130_fd_sc_hd__nand2_1 _10284_ (.A(_02517_),
    .B(_02518_),
    .Y(_02519_));
 sky130_fd_sc_hd__and4_1 _10285_ (.A(_02159_),
    .B(_02505_),
    .C(_02506_),
    .D(_02519_),
    .X(_02520_));
 sky130_fd_sc_hd__a31o_1 _10286_ (.A1(_02159_),
    .A2(_02505_),
    .A3(_02506_),
    .B1(_02519_),
    .X(_02522_));
 sky130_fd_sc_hd__and2b_1 _10287_ (.A_N(_02520_),
    .B(_02522_),
    .X(_02523_));
 sky130_fd_sc_hd__and3_1 _10288_ (.A(_00628_),
    .B(_05742_),
    .C(_01545_),
    .X(_02524_));
 sky130_fd_sc_hd__a22o_1 _10289_ (.A1(_05742_),
    .A2(_01545_),
    .B1(_02156_),
    .B2(_00628_),
    .X(_02525_));
 sky130_fd_sc_hd__a21bo_1 _10290_ (.A1(_02156_),
    .A2(_02524_),
    .B1_N(_02525_),
    .X(_02526_));
 sky130_fd_sc_hd__nand2_1 _10291_ (.A(_05577_),
    .B(_01410_),
    .Y(_02527_));
 sky130_fd_sc_hd__xor2_1 _10292_ (.A(_02526_),
    .B(_02527_),
    .X(_02528_));
 sky130_fd_sc_hd__a31o_1 _10293_ (.A1(_05577_),
    .A2(net49),
    .A3(_02326_),
    .B1(_02323_),
    .X(_02529_));
 sky130_fd_sc_hd__nand2_1 _10294_ (.A(_03268_),
    .B(_01058_),
    .Y(_02530_));
 sky130_fd_sc_hd__xnor2_1 _10295_ (.A(_02529_),
    .B(_02530_),
    .Y(_02531_));
 sky130_fd_sc_hd__xor2_1 _10296_ (.A(_02528_),
    .B(_02531_),
    .X(_02533_));
 sky130_fd_sc_hd__nand2_1 _10297_ (.A(_02329_),
    .B(_02533_),
    .Y(_02534_));
 sky130_fd_sc_hd__or2_1 _10298_ (.A(_02329_),
    .B(_02533_),
    .X(_02535_));
 sky130_fd_sc_hd__nand2_1 _10299_ (.A(_02534_),
    .B(_02535_),
    .Y(_02536_));
 sky130_fd_sc_hd__xnor2_2 _10300_ (.A(_02523_),
    .B(_02536_),
    .Y(_02537_));
 sky130_fd_sc_hd__xnor2_2 _10301_ (.A(_02504_),
    .B(_02537_),
    .Y(_02538_));
 sky130_fd_sc_hd__nand2_1 _10302_ (.A(_02301_),
    .B(_02332_),
    .Y(_02539_));
 sky130_fd_sc_hd__o21ai_2 _10303_ (.A1(_02180_),
    .A2(_02333_),
    .B1(_02539_),
    .Y(_02540_));
 sky130_fd_sc_hd__xor2_2 _10304_ (.A(_02538_),
    .B(_02540_),
    .X(_02541_));
 sky130_fd_sc_hd__xnor2_1 _10305_ (.A(_02502_),
    .B(_02541_),
    .Y(_02542_));
 sky130_fd_sc_hd__o21ba_1 _10306_ (.A1(_02355_),
    .A2(_02363_),
    .B1_N(_02374_),
    .X(_02544_));
 sky130_fd_sc_hd__a21o_2 _10307_ (.A1(_02355_),
    .A2(_02363_),
    .B1(_02544_),
    .X(_02545_));
 sky130_fd_sc_hd__nand2_1 _10308_ (.A(_02350_),
    .B(_02352_),
    .Y(_02546_));
 sky130_fd_sc_hd__nand2_1 _10309_ (.A(_02353_),
    .B(_02354_),
    .Y(_02547_));
 sky130_fd_sc_hd__and3_1 _10310_ (.A(_00366_),
    .B(_02971_),
    .C(_01368_),
    .X(_02548_));
 sky130_fd_sc_hd__a22o_1 _10311_ (.A1(_02971_),
    .A2(_01368_),
    .B1(_00959_),
    .B2(_00366_),
    .X(_02549_));
 sky130_fd_sc_hd__a21bo_1 _10312_ (.A1(_01369_),
    .A2(_02548_),
    .B1_N(_02549_),
    .X(_02550_));
 sky130_fd_sc_hd__nand2_1 _10313_ (.A(_05203_),
    .B(_00604_),
    .Y(_02551_));
 sky130_fd_sc_hd__xor2_1 _10314_ (.A(_02550_),
    .B(_02551_),
    .X(_02552_));
 sky130_fd_sc_hd__a32o_1 _10315_ (.A1(_05192_),
    .A2(net45),
    .A3(_02356_),
    .B1(_02224_),
    .B2(_01506_),
    .X(_02553_));
 sky130_fd_sc_hd__nand2_1 _10316_ (.A(_04598_),
    .B(net45),
    .Y(_02555_));
 sky130_fd_sc_hd__xnor2_1 _10317_ (.A(_02553_),
    .B(_02555_),
    .Y(_02556_));
 sky130_fd_sc_hd__xor2_1 _10318_ (.A(_02552_),
    .B(_02556_),
    .X(_02557_));
 sky130_fd_sc_hd__nand2_1 _10319_ (.A(_02361_),
    .B(_02557_),
    .Y(_02558_));
 sky130_fd_sc_hd__or2_1 _10320_ (.A(_02361_),
    .B(_02557_),
    .X(_02559_));
 sky130_fd_sc_hd__nand2_1 _10321_ (.A(_02558_),
    .B(_02559_),
    .Y(_02560_));
 sky130_fd_sc_hd__and4_1 _10322_ (.A(_02214_),
    .B(_02546_),
    .C(_02547_),
    .D(_02560_),
    .X(_02561_));
 sky130_fd_sc_hd__a31o_1 _10323_ (.A1(_02214_),
    .A2(_02546_),
    .A3(_02547_),
    .B1(_02560_),
    .X(_02562_));
 sky130_fd_sc_hd__and2b_1 _10324_ (.A_N(_02561_),
    .B(_02562_),
    .X(_02563_));
 sky130_fd_sc_hd__and3_1 _10325_ (.A(_04862_),
    .B(net4),
    .C(_00780_),
    .X(_02564_));
 sky130_fd_sc_hd__a22o_1 _10326_ (.A1(_04851_),
    .A2(_00780_),
    .B1(_00777_),
    .B2(net4),
    .X(_02566_));
 sky130_fd_sc_hd__a21bo_1 _10327_ (.A1(_00613_),
    .A2(_02564_),
    .B1_N(_02566_),
    .X(_02567_));
 sky130_fd_sc_hd__nand2_1 _10328_ (.A(_05027_),
    .B(_00373_),
    .Y(_02568_));
 sky130_fd_sc_hd__xor2_1 _10329_ (.A(_02567_),
    .B(_02568_),
    .X(_02569_));
 sky130_fd_sc_hd__a31o_1 _10330_ (.A1(_05027_),
    .A2(net40),
    .A3(_02369_),
    .B1(_02366_),
    .X(_02570_));
 sky130_fd_sc_hd__nand2_1 _10331_ (.A(net7),
    .B(_04048_),
    .Y(_02571_));
 sky130_fd_sc_hd__xnor2_1 _10332_ (.A(_02570_),
    .B(_02571_),
    .Y(_02572_));
 sky130_fd_sc_hd__xor2_1 _10333_ (.A(_02569_),
    .B(_02572_),
    .X(_02573_));
 sky130_fd_sc_hd__nand2_1 _10334_ (.A(_02372_),
    .B(_02573_),
    .Y(_02574_));
 sky130_fd_sc_hd__or2_1 _10335_ (.A(_02372_),
    .B(_02573_),
    .X(_02575_));
 sky130_fd_sc_hd__nand2_2 _10336_ (.A(_02574_),
    .B(_02575_),
    .Y(_02577_));
 sky130_fd_sc_hd__xnor2_4 _10337_ (.A(_02563_),
    .B(_02577_),
    .Y(_02578_));
 sky130_fd_sc_hd__xor2_4 _10338_ (.A(_02545_),
    .B(_02578_),
    .X(_02579_));
 sky130_fd_sc_hd__nand2_1 _10339_ (.A(_02349_),
    .B(_02375_),
    .Y(_02580_));
 sky130_fd_sc_hd__o21ai_4 _10340_ (.A1(_02233_),
    .A2(_02376_),
    .B1(_02580_),
    .Y(_02581_));
 sky130_fd_sc_hd__xnor2_4 _10341_ (.A(_02579_),
    .B(_02581_),
    .Y(_02582_));
 sky130_fd_sc_hd__xnor2_2 _10342_ (.A(_02542_),
    .B(_02582_),
    .Y(_02583_));
 sky130_fd_sc_hd__nand2_1 _10343_ (.A(_02334_),
    .B(_02345_),
    .Y(_02584_));
 sky130_fd_sc_hd__nor2_1 _10344_ (.A(_02334_),
    .B(_02345_),
    .Y(_02585_));
 sky130_fd_sc_hd__a21oi_2 _10345_ (.A1(_02584_),
    .A2(_02377_),
    .B1(_02585_),
    .Y(_02586_));
 sky130_fd_sc_hd__xnor2_2 _10346_ (.A(_02583_),
    .B(_02586_),
    .Y(_02588_));
 sky130_fd_sc_hd__a21o_1 _10347_ (.A1(_02382_),
    .A2(_02385_),
    .B1(_02588_),
    .X(_02589_));
 sky130_fd_sc_hd__nand3_1 _10348_ (.A(_02382_),
    .B(_02385_),
    .C(_02588_),
    .Y(_02590_));
 sky130_fd_sc_hd__nand2_1 _10349_ (.A(_02589_),
    .B(_02590_),
    .Y(_02591_));
 sky130_fd_sc_hd__a21o_1 _10350_ (.A1(_02496_),
    .A2(_02498_),
    .B1(_02591_),
    .X(_02592_));
 sky130_fd_sc_hd__nand3_1 _10351_ (.A(_02496_),
    .B(_02498_),
    .C(_02591_),
    .Y(_02593_));
 sky130_fd_sc_hd__inv_2 _10352_ (.A(_02433_),
    .Y(_02594_));
 sky130_fd_sc_hd__a211oi_1 _10353_ (.A1(_02095_),
    .A2(_02429_),
    .B1(_02432_),
    .C1(_02092_),
    .Y(_02595_));
 sky130_fd_sc_hd__o21ai_2 _10354_ (.A1(_02594_),
    .A2(_02436_),
    .B1(_02595_),
    .Y(_02596_));
 sky130_fd_sc_hd__inv_2 _10355_ (.A(_02065_),
    .Y(_02597_));
 sky130_fd_sc_hd__and2_1 _10356_ (.A(_02397_),
    .B(_02398_),
    .X(_02599_));
 sky130_fd_sc_hd__and3_1 _10357_ (.A(_07010_),
    .B(_00101_),
    .C(_00423_),
    .X(_02600_));
 sky130_fd_sc_hd__a22o_1 _10358_ (.A1(_07010_),
    .A2(_03685_),
    .B1(_00423_),
    .B2(_00101_),
    .X(_02601_));
 sky130_fd_sc_hd__a21bo_1 _10359_ (.A1(_03696_),
    .A2(_02600_),
    .B1_N(_02601_),
    .X(_02602_));
 sky130_fd_sc_hd__nand2_1 _10360_ (.A(_06733_),
    .B(_03773_),
    .Y(_02603_));
 sky130_fd_sc_hd__xor2_1 _10361_ (.A(_02602_),
    .B(_02603_),
    .X(_02604_));
 sky130_fd_sc_hd__a31o_1 _10362_ (.A1(_06744_),
    .A2(_03894_),
    .A3(_02400_),
    .B1(_02403_),
    .X(_02605_));
 sky130_fd_sc_hd__nand2_1 _10363_ (.A(_06744_),
    .B(_03938_),
    .Y(_02606_));
 sky130_fd_sc_hd__xnor2_1 _10364_ (.A(_02605_),
    .B(_02606_),
    .Y(_02607_));
 sky130_fd_sc_hd__nand2_1 _10365_ (.A(_02604_),
    .B(_02607_),
    .Y(_02608_));
 sky130_fd_sc_hd__or2_1 _10366_ (.A(_02604_),
    .B(_02607_),
    .X(_02610_));
 sky130_fd_sc_hd__nand2_1 _10367_ (.A(_02608_),
    .B(_02610_),
    .Y(_02611_));
 sky130_fd_sc_hd__nor2_1 _10368_ (.A(_02407_),
    .B(_02611_),
    .Y(_02612_));
 sky130_fd_sc_hd__and2_1 _10369_ (.A(_02407_),
    .B(_02611_),
    .X(_02613_));
 sky130_fd_sc_hd__nor2_1 _10370_ (.A(_02612_),
    .B(_02613_),
    .Y(_02614_));
 sky130_fd_sc_hd__or4_2 _10371_ (.A(_02597_),
    .B(_02395_),
    .C(_02599_),
    .D(_02614_),
    .X(_02615_));
 sky130_fd_sc_hd__o31ai_2 _10372_ (.A1(_02597_),
    .A2(_02395_),
    .A3(_02599_),
    .B1(_02614_),
    .Y(_02616_));
 sky130_fd_sc_hd__nand2_1 _10373_ (.A(_02615_),
    .B(_02616_),
    .Y(_02617_));
 sky130_fd_sc_hd__and3_1 _10374_ (.A(_06819_),
    .B(_06821_),
    .C(_00730_),
    .X(_02618_));
 sky130_fd_sc_hd__a22o_1 _10375_ (.A1(_06819_),
    .A2(_00413_),
    .B1(_00571_),
    .B2(_06821_),
    .X(_02619_));
 sky130_fd_sc_hd__a21bo_1 _10376_ (.A1(_00413_),
    .A2(_02618_),
    .B1_N(_02619_),
    .X(_02621_));
 sky130_fd_sc_hd__nand2_1 _10377_ (.A(_03521_),
    .B(_00734_),
    .Y(_02622_));
 sky130_fd_sc_hd__xor2_1 _10378_ (.A(_02621_),
    .B(_02622_),
    .X(_02623_));
 sky130_fd_sc_hd__a31o_1 _10379_ (.A1(_00475_),
    .A2(_00734_),
    .A3(_02411_),
    .B1(_02414_),
    .X(_02624_));
 sky130_fd_sc_hd__nand2_1 _10380_ (.A(_00486_),
    .B(_01211_),
    .Y(_02625_));
 sky130_fd_sc_hd__xnor2_1 _10381_ (.A(_02624_),
    .B(_02625_),
    .Y(_02626_));
 sky130_fd_sc_hd__nand2_1 _10382_ (.A(_02623_),
    .B(_02626_),
    .Y(_02627_));
 sky130_fd_sc_hd__or2_1 _10383_ (.A(_02623_),
    .B(_02626_),
    .X(_02628_));
 sky130_fd_sc_hd__nand2_1 _10384_ (.A(_02627_),
    .B(_02628_),
    .Y(_02629_));
 sky130_fd_sc_hd__nor2_1 _10385_ (.A(_02418_),
    .B(_02629_),
    .Y(_02630_));
 sky130_fd_sc_hd__and2_1 _10386_ (.A(_02418_),
    .B(_02629_),
    .X(_02632_));
 sky130_fd_sc_hd__or2_1 _10387_ (.A(_02630_),
    .B(_02632_),
    .X(_02633_));
 sky130_fd_sc_hd__xor2_1 _10388_ (.A(_02617_),
    .B(_02633_),
    .X(_02634_));
 sky130_fd_sc_hd__nand2_1 _10389_ (.A(_02399_),
    .B(_02409_),
    .Y(_02635_));
 sky130_fd_sc_hd__o21ai_1 _10390_ (.A1(_02399_),
    .A2(_02409_),
    .B1(_02420_),
    .Y(_02636_));
 sky130_fd_sc_hd__nand2_1 _10391_ (.A(_02635_),
    .B(_02636_),
    .Y(_02637_));
 sky130_fd_sc_hd__and2b_1 _10392_ (.A_N(_02634_),
    .B(_02637_),
    .X(_02638_));
 sky130_fd_sc_hd__and3_1 _10393_ (.A(_02635_),
    .B(_02636_),
    .C(_02634_),
    .X(_02639_));
 sky130_fd_sc_hd__or2_1 _10394_ (.A(_02638_),
    .B(_02639_),
    .X(_02640_));
 sky130_fd_sc_hd__and2_1 _10395_ (.A(_02392_),
    .B(_02421_),
    .X(_02641_));
 sky130_fd_sc_hd__a21o_1 _10396_ (.A1(_02082_),
    .A2(_02422_),
    .B1(_02641_),
    .X(_02643_));
 sky130_fd_sc_hd__xnor2_2 _10397_ (.A(_02640_),
    .B(_02643_),
    .Y(_02644_));
 sky130_fd_sc_hd__xnor2_1 _10398_ (.A(_02596_),
    .B(_02644_),
    .Y(_02645_));
 sky130_fd_sc_hd__inv_2 _10399_ (.A(_02121_),
    .Y(_02646_));
 sky130_fd_sc_hd__and2_1 _10400_ (.A(_02444_),
    .B(_02446_),
    .X(_02647_));
 sky130_fd_sc_hd__and3_1 _10401_ (.A(_05445_),
    .B(_05467_),
    .C(_01246_),
    .X(_02648_));
 sky130_fd_sc_hd__a22o_1 _10402_ (.A1(_05445_),
    .A2(_01177_),
    .B1(_01247_),
    .B2(_05467_),
    .X(_02649_));
 sky130_fd_sc_hd__a21bo_1 _10403_ (.A1(_01178_),
    .A2(_02648_),
    .B1_N(_02649_),
    .X(_02650_));
 sky130_fd_sc_hd__nand2_1 _10404_ (.A(_02007_),
    .B(_02117_),
    .Y(_02651_));
 sky130_fd_sc_hd__xor2_1 _10405_ (.A(_02650_),
    .B(_02651_),
    .X(_02652_));
 sky130_fd_sc_hd__a31o_1 _10406_ (.A1(_02029_),
    .A2(_01564_),
    .A3(_02448_),
    .B1(_02450_),
    .X(_02654_));
 sky130_fd_sc_hd__nand2_1 _10407_ (.A(_02029_),
    .B(_01960_),
    .Y(_02655_));
 sky130_fd_sc_hd__xnor2_1 _10408_ (.A(_02654_),
    .B(_02655_),
    .Y(_02656_));
 sky130_fd_sc_hd__nand2_1 _10409_ (.A(_02652_),
    .B(_02656_),
    .Y(_02657_));
 sky130_fd_sc_hd__or2_1 _10410_ (.A(_02652_),
    .B(_02656_),
    .X(_02658_));
 sky130_fd_sc_hd__nand2_1 _10411_ (.A(_02657_),
    .B(_02658_),
    .Y(_02659_));
 sky130_fd_sc_hd__nor2_1 _10412_ (.A(_02454_),
    .B(_02659_),
    .Y(_02660_));
 sky130_fd_sc_hd__and2_1 _10413_ (.A(_02454_),
    .B(_02659_),
    .X(_02661_));
 sky130_fd_sc_hd__nor2_1 _10414_ (.A(_02660_),
    .B(_02661_),
    .Y(_02662_));
 sky130_fd_sc_hd__or4_2 _10415_ (.A(_02646_),
    .B(_02442_),
    .C(_02647_),
    .D(_02662_),
    .X(_02663_));
 sky130_fd_sc_hd__o31ai_2 _10416_ (.A1(_02646_),
    .A2(_02442_),
    .A3(_02647_),
    .B1(_02662_),
    .Y(_02665_));
 sky130_fd_sc_hd__nand2_1 _10417_ (.A(_02663_),
    .B(_02665_),
    .Y(_02666_));
 sky130_fd_sc_hd__and3_1 _10418_ (.A(_01295_),
    .B(_01306_),
    .C(net22),
    .X(_02667_));
 sky130_fd_sc_hd__a22o_1 _10419_ (.A1(_01295_),
    .A2(net21),
    .B1(_02133_),
    .B2(_01306_),
    .X(_02668_));
 sky130_fd_sc_hd__a21bo_1 _10420_ (.A1(net21),
    .A2(_02667_),
    .B1_N(_02668_),
    .X(_02669_));
 sky130_fd_sc_hd__nand2_1 _10421_ (.A(_02127_),
    .B(_02459_),
    .Y(_02670_));
 sky130_fd_sc_hd__xor2_1 _10422_ (.A(_02669_),
    .B(_02670_),
    .X(_02671_));
 sky130_fd_sc_hd__a31o_1 _10423_ (.A1(_00311_),
    .A2(net24),
    .A3(_02460_),
    .B1(_02462_),
    .X(_02672_));
 sky130_fd_sc_hd__clkbuf_4 _10424_ (.A(net25),
    .X(_02673_));
 sky130_fd_sc_hd__nand2_1 _10425_ (.A(_00322_),
    .B(_02673_),
    .Y(_02674_));
 sky130_fd_sc_hd__xnor2_1 _10426_ (.A(_02672_),
    .B(_02674_),
    .Y(_02676_));
 sky130_fd_sc_hd__nand2_1 _10427_ (.A(_02671_),
    .B(_02676_),
    .Y(_02677_));
 sky130_fd_sc_hd__or2_1 _10428_ (.A(_02671_),
    .B(_02676_),
    .X(_02678_));
 sky130_fd_sc_hd__nand2_1 _10429_ (.A(_02677_),
    .B(_02678_),
    .Y(_02679_));
 sky130_fd_sc_hd__nor2_1 _10430_ (.A(_02466_),
    .B(_02679_),
    .Y(_02680_));
 sky130_fd_sc_hd__and2_1 _10431_ (.A(_02466_),
    .B(_02679_),
    .X(_02681_));
 sky130_fd_sc_hd__or2_1 _10432_ (.A(_02680_),
    .B(_02681_),
    .X(_02682_));
 sky130_fd_sc_hd__xor2_1 _10433_ (.A(_02666_),
    .B(_02682_),
    .X(_02683_));
 sky130_fd_sc_hd__nand2_1 _10434_ (.A(_02447_),
    .B(_02457_),
    .Y(_02684_));
 sky130_fd_sc_hd__o21ai_1 _10435_ (.A1(_02447_),
    .A2(_02457_),
    .B1(_02469_),
    .Y(_02685_));
 sky130_fd_sc_hd__nand2_1 _10436_ (.A(_02684_),
    .B(_02685_),
    .Y(_02687_));
 sky130_fd_sc_hd__and2b_1 _10437_ (.A_N(_02683_),
    .B(_02687_),
    .X(_02688_));
 sky130_fd_sc_hd__and3_1 _10438_ (.A(_02684_),
    .B(_02685_),
    .C(_02683_),
    .X(_02689_));
 sky130_fd_sc_hd__or2_2 _10439_ (.A(_02688_),
    .B(_02689_),
    .X(_02690_));
 sky130_fd_sc_hd__and2_1 _10440_ (.A(_02439_),
    .B(_02470_),
    .X(_02691_));
 sky130_fd_sc_hd__a21o_2 _10441_ (.A1(_02142_),
    .A2(_02471_),
    .B1(_02691_),
    .X(_02692_));
 sky130_fd_sc_hd__xnor2_4 _10442_ (.A(_02690_),
    .B(_02692_),
    .Y(_02693_));
 sky130_fd_sc_hd__xnor2_2 _10443_ (.A(_02645_),
    .B(_02693_),
    .Y(_02694_));
 sky130_fd_sc_hd__nand2_1 _10444_ (.A(_02424_),
    .B(_02437_),
    .Y(_02695_));
 sky130_fd_sc_hd__nor2_1 _10445_ (.A(_02424_),
    .B(_02437_),
    .Y(_02696_));
 sky130_fd_sc_hd__a21oi_2 _10446_ (.A1(_02695_),
    .A2(_02472_),
    .B1(_02696_),
    .Y(_02698_));
 sky130_fd_sc_hd__xnor2_2 _10447_ (.A(_02694_),
    .B(_02698_),
    .Y(_02699_));
 sky130_fd_sc_hd__nor2_1 _10448_ (.A(_02476_),
    .B(_02480_),
    .Y(_02700_));
 sky130_fd_sc_hd__or2_2 _10449_ (.A(_02699_),
    .B(_02700_),
    .X(_02701_));
 sky130_fd_sc_hd__nand2_1 _10450_ (.A(_02699_),
    .B(_02700_),
    .Y(_02702_));
 sky130_fd_sc_hd__nand2_4 _10451_ (.A(_02701_),
    .B(_02702_),
    .Y(_02703_));
 sky130_fd_sc_hd__nand3_1 _10452_ (.A(_02592_),
    .B(_02593_),
    .C(_02703_),
    .Y(_02704_));
 sky130_fd_sc_hd__a21o_1 _10453_ (.A1(_02592_),
    .A2(_02593_),
    .B1(_02703_),
    .X(_02705_));
 sky130_fd_sc_hd__inv_2 _10454_ (.A(_02482_),
    .Y(_02706_));
 sky130_fd_sc_hd__a21boi_2 _10455_ (.A1(_02389_),
    .A2(_02706_),
    .B1_N(_02388_),
    .Y(_02707_));
 sky130_fd_sc_hd__a21o_2 _10456_ (.A1(_02704_),
    .A2(_02705_),
    .B1(_02707_),
    .X(_02709_));
 sky130_fd_sc_hd__nand3_1 _10457_ (.A(_02704_),
    .B(_02705_),
    .C(_02707_),
    .Y(_02710_));
 sky130_fd_sc_hd__and3_1 _10458_ (.A(_02487_),
    .B(_02709_),
    .C(_02710_),
    .X(_02711_));
 sky130_fd_sc_hd__a21oi_1 _10459_ (.A1(_02709_),
    .A2(_02710_),
    .B1(_02487_),
    .Y(_02712_));
 sky130_fd_sc_hd__nor2_4 _10460_ (.A(_02711_),
    .B(_02712_),
    .Y(_02713_));
 sky130_fd_sc_hd__and2_1 _10461_ (.A(_02274_),
    .B(_02491_),
    .X(_02714_));
 sky130_fd_sc_hd__a21o_1 _10462_ (.A1(_02052_),
    .A2(_02273_),
    .B1(_02279_),
    .X(_02715_));
 sky130_fd_sc_hd__inv_2 _10463_ (.A(_02490_),
    .Y(_02716_));
 sky130_fd_sc_hd__a32o_1 _10464_ (.A1(_02274_),
    .A2(_02276_),
    .A3(_02491_),
    .B1(_02715_),
    .B2(_02716_),
    .X(_02717_));
 sky130_fd_sc_hd__a31o_1 _10465_ (.A1(_01649_),
    .A2(_02275_),
    .A3(_02714_),
    .B1(_02717_),
    .X(_02718_));
 sky130_fd_sc_hd__xor2_4 _10466_ (.A(_02713_),
    .B(_02718_),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_4 _10467_ (.A(_02169_),
    .X(_02720_));
 sky130_fd_sc_hd__clkbuf_4 _10468_ (.A(_02720_),
    .X(_02721_));
 sky130_fd_sc_hd__clkbuf_4 _10469_ (.A(_02721_),
    .X(_02722_));
 sky130_fd_sc_hd__buf_2 _10470_ (.A(_02312_),
    .X(_02723_));
 sky130_fd_sc_hd__clkbuf_4 _10471_ (.A(_02723_),
    .X(_02724_));
 sky130_fd_sc_hd__clkbuf_4 _10472_ (.A(_02724_),
    .X(_02725_));
 sky130_fd_sc_hd__clkbuf_4 _10473_ (.A(_02725_),
    .X(_02726_));
 sky130_fd_sc_hd__clkbuf_4 _10474_ (.A(net57),
    .X(_02727_));
 sky130_fd_sc_hd__clkbuf_4 _10475_ (.A(_02727_),
    .X(_02728_));
 sky130_fd_sc_hd__clkbuf_4 _10476_ (.A(_02728_),
    .X(_02730_));
 sky130_fd_sc_hd__clkbuf_4 _10477_ (.A(_02730_),
    .X(_02731_));
 sky130_fd_sc_hd__a22o_1 _10478_ (.A1(_01472_),
    .A2(_02726_),
    .B1(_02731_),
    .B2(_00636_),
    .X(_02732_));
 sky130_fd_sc_hd__and4_1 _10479_ (.A(_01472_),
    .B(_00636_),
    .C(_02726_),
    .D(_02730_),
    .X(_02733_));
 sky130_fd_sc_hd__a31o_1 _10480_ (.A1(_02247_),
    .A2(_02722_),
    .A3(_02732_),
    .B1(_02733_),
    .X(_02734_));
 sky130_fd_sc_hd__clkbuf_4 _10481_ (.A(_02726_),
    .X(_02735_));
 sky130_fd_sc_hd__clkbuf_4 _10482_ (.A(_02735_),
    .X(_02736_));
 sky130_fd_sc_hd__clkbuf_4 _10483_ (.A(_02731_),
    .X(_02737_));
 sky130_fd_sc_hd__nand4_1 _10484_ (.A(_01473_),
    .B(_02247_),
    .C(_02736_),
    .D(_02737_),
    .Y(_02738_));
 sky130_fd_sc_hd__a22o_1 _10485_ (.A1(_02247_),
    .A2(_02736_),
    .B1(_02737_),
    .B2(_01473_),
    .X(_02739_));
 sky130_fd_sc_hd__and3_1 _10486_ (.A(_02734_),
    .B(_02738_),
    .C(_02739_),
    .X(_02741_));
 sky130_fd_sc_hd__clkbuf_4 _10487_ (.A(_02737_),
    .X(_02742_));
 sky130_fd_sc_hd__clkbuf_4 _10488_ (.A(_02736_),
    .X(_02743_));
 sky130_fd_sc_hd__nand2_1 _10489_ (.A(_01473_),
    .B(_02743_),
    .Y(_02744_));
 sky130_fd_sc_hd__and3_1 _10490_ (.A(_02247_),
    .B(_02742_),
    .C(_02744_),
    .X(_02745_));
 sky130_fd_sc_hd__xor2_2 _10491_ (.A(_02741_),
    .B(_02745_),
    .X(_02746_));
 sky130_fd_sc_hd__or2b_1 _10492_ (.A(_02733_),
    .B_N(_02732_),
    .X(_02747_));
 sky130_fd_sc_hd__nand2_1 _10493_ (.A(_02247_),
    .B(_02721_),
    .Y(_02748_));
 sky130_fd_sc_hd__xnor2_1 _10494_ (.A(_02747_),
    .B(_02748_),
    .Y(_02749_));
 sky130_fd_sc_hd__a22o_1 _10495_ (.A1(_00636_),
    .A2(_02735_),
    .B1(_02731_),
    .B2(_00526_),
    .X(_02750_));
 sky130_fd_sc_hd__and4_1 _10496_ (.A(_00636_),
    .B(_00526_),
    .C(_02735_),
    .D(_02731_),
    .X(_02752_));
 sky130_fd_sc_hd__a31o_1 _10497_ (.A1(_01473_),
    .A2(_02721_),
    .A3(_02750_),
    .B1(_02752_),
    .X(_02753_));
 sky130_fd_sc_hd__and2b_1 _10498_ (.A_N(_02749_),
    .B(_02753_),
    .X(_02754_));
 sky130_fd_sc_hd__a21oi_1 _10499_ (.A1(_02738_),
    .A2(_02739_),
    .B1(_02734_),
    .Y(_02755_));
 sky130_fd_sc_hd__nor2_1 _10500_ (.A(_02741_),
    .B(_02755_),
    .Y(_02756_));
 sky130_fd_sc_hd__xnor2_1 _10501_ (.A(_02754_),
    .B(_02756_),
    .Y(_02757_));
 sky130_fd_sc_hd__clkbuf_4 _10502_ (.A(_01934_),
    .X(_02758_));
 sky130_fd_sc_hd__clkbuf_4 _10503_ (.A(_02758_),
    .X(_02759_));
 sky130_fd_sc_hd__and4_1 _10504_ (.A(_00635_),
    .B(_07040_),
    .C(_02720_),
    .D(_02726_),
    .X(_02760_));
 sky130_fd_sc_hd__inv_2 _10505_ (.A(_02760_),
    .Y(_02761_));
 sky130_fd_sc_hd__a22o_1 _10506_ (.A1(_00636_),
    .A2(_02721_),
    .B1(_02726_),
    .B2(_00526_),
    .X(_02763_));
 sky130_fd_sc_hd__and4_1 _10507_ (.A(_01472_),
    .B(_02759_),
    .C(_02761_),
    .D(_02763_),
    .X(_02764_));
 sky130_fd_sc_hd__clkbuf_4 _10508_ (.A(_02759_),
    .X(_02765_));
 sky130_fd_sc_hd__clkbuf_4 _10509_ (.A(_02765_),
    .X(_02766_));
 sky130_fd_sc_hd__a22oi_1 _10510_ (.A1(_01473_),
    .A2(_02766_),
    .B1(_02761_),
    .B2(_02763_),
    .Y(_02767_));
 sky130_fd_sc_hd__nor2_1 _10511_ (.A(_02764_),
    .B(_02767_),
    .Y(_02768_));
 sky130_fd_sc_hd__and4_1 _10512_ (.A(_00636_),
    .B(_01156_),
    .C(_02765_),
    .D(_02722_),
    .X(_02769_));
 sky130_fd_sc_hd__nand2_1 _10513_ (.A(_02768_),
    .B(_02769_),
    .Y(_02770_));
 sky130_fd_sc_hd__nand2_1 _10514_ (.A(_02247_),
    .B(_02765_),
    .Y(_02771_));
 sky130_fd_sc_hd__or2_1 _10515_ (.A(_02760_),
    .B(_02764_),
    .X(_02772_));
 sky130_fd_sc_hd__or2b_1 _10516_ (.A(_02771_),
    .B_N(_02772_),
    .X(_02774_));
 sky130_fd_sc_hd__and2b_1 _10517_ (.A_N(_02752_),
    .B(_02750_),
    .X(_02775_));
 sky130_fd_sc_hd__nand2_1 _10518_ (.A(_01473_),
    .B(_02722_),
    .Y(_02776_));
 sky130_fd_sc_hd__xnor2_1 _10519_ (.A(_02775_),
    .B(_02776_),
    .Y(_02777_));
 sky130_fd_sc_hd__xnor2_1 _10520_ (.A(_02772_),
    .B(_02771_),
    .Y(_02778_));
 sky130_fd_sc_hd__nand2_1 _10521_ (.A(_02777_),
    .B(_02778_),
    .Y(_02779_));
 sky130_fd_sc_hd__and2b_1 _10522_ (.A_N(_02753_),
    .B(_02749_),
    .X(_02780_));
 sky130_fd_sc_hd__or2_1 _10523_ (.A(_02754_),
    .B(_02780_),
    .X(_02781_));
 sky130_fd_sc_hd__a21o_1 _10524_ (.A1(_02774_),
    .A2(_02779_),
    .B1(_02781_),
    .X(_02782_));
 sky130_fd_sc_hd__nand3_1 _10525_ (.A(_02774_),
    .B(_02779_),
    .C(_02781_),
    .Y(_02783_));
 sky130_fd_sc_hd__nand2_1 _10526_ (.A(_02782_),
    .B(_02783_),
    .Y(_02785_));
 sky130_fd_sc_hd__or2_1 _10527_ (.A(_02777_),
    .B(_02778_),
    .X(_02786_));
 sky130_fd_sc_hd__nand2_1 _10528_ (.A(_02779_),
    .B(_02786_),
    .Y(_02787_));
 sky130_fd_sc_hd__o31a_1 _10529_ (.A1(_02770_),
    .A2(_02785_),
    .A3(_02787_),
    .B1(_02782_),
    .X(_02788_));
 sky130_fd_sc_hd__nor2_1 _10530_ (.A(_02757_),
    .B(_02788_),
    .Y(_02789_));
 sky130_fd_sc_hd__a21o_1 _10531_ (.A1(_02754_),
    .A2(_02756_),
    .B1(_02789_),
    .X(_02790_));
 sky130_fd_sc_hd__a21bo_1 _10532_ (.A1(_02741_),
    .A2(_02745_),
    .B1_N(_02738_),
    .X(_02791_));
 sky130_fd_sc_hd__a21oi_1 _10533_ (.A1(_02746_),
    .A2(_02790_),
    .B1(_02791_),
    .Y(_02792_));
 sky130_fd_sc_hd__inv_2 _10534_ (.A(_02792_),
    .Y(_02793_));
 sky130_fd_sc_hd__or2_1 _10535_ (.A(_02768_),
    .B(_02769_),
    .X(_02794_));
 sky130_fd_sc_hd__nand2_2 _10536_ (.A(_02770_),
    .B(_02794_),
    .Y(_02796_));
 sky130_fd_sc_hd__and4_1 _10537_ (.A(_03004_),
    .B(_00293_),
    .C(_02724_),
    .D(_02728_),
    .X(_02797_));
 sky130_fd_sc_hd__a22o_1 _10538_ (.A1(_00293_),
    .A2(_02725_),
    .B1(_02728_),
    .B2(_03015_),
    .X(_02798_));
 sky130_fd_sc_hd__or2b_1 _10539_ (.A(_02797_),
    .B_N(_02798_),
    .X(_02799_));
 sky130_fd_sc_hd__nand2_1 _10540_ (.A(_00294_),
    .B(_02169_),
    .Y(_02800_));
 sky130_fd_sc_hd__xnor2_1 _10541_ (.A(_02799_),
    .B(_02800_),
    .Y(_02801_));
 sky130_fd_sc_hd__a22o_1 _10542_ (.A1(_03004_),
    .A2(_02724_),
    .B1(_02728_),
    .B2(_00388_),
    .X(_02802_));
 sky130_fd_sc_hd__and4_1 _10543_ (.A(_00388_),
    .B(_03004_),
    .C(_02724_),
    .D(_02727_),
    .X(_02803_));
 sky130_fd_sc_hd__a31o_1 _10544_ (.A1(_00819_),
    .A2(_02169_),
    .A3(_02802_),
    .B1(_02803_),
    .X(_02804_));
 sky130_fd_sc_hd__or2b_1 _10545_ (.A(_02801_),
    .B_N(_02804_),
    .X(_02805_));
 sky130_fd_sc_hd__a31o_1 _10546_ (.A1(_00818_),
    .A2(_02169_),
    .A3(_02798_),
    .B1(_02797_),
    .X(_02807_));
 sky130_fd_sc_hd__nand4_1 _10547_ (.A(_00819_),
    .B(_00818_),
    .C(_02725_),
    .D(_02730_),
    .Y(_02808_));
 sky130_fd_sc_hd__a22o_1 _10548_ (.A1(_00818_),
    .A2(_02725_),
    .B1(_02730_),
    .B2(_00819_),
    .X(_02809_));
 sky130_fd_sc_hd__and3_1 _10549_ (.A(_02807_),
    .B(_02808_),
    .C(_02809_),
    .X(_02810_));
 sky130_fd_sc_hd__a21oi_1 _10550_ (.A1(_02808_),
    .A2(_02809_),
    .B1(_02807_),
    .Y(_02811_));
 sky130_fd_sc_hd__nor2_1 _10551_ (.A(_02810_),
    .B(_02811_),
    .Y(_02812_));
 sky130_fd_sc_hd__xor2_1 _10552_ (.A(_02805_),
    .B(_02812_),
    .X(_02813_));
 sky130_fd_sc_hd__and4_1 _10553_ (.A(_00377_),
    .B(_02993_),
    .C(_02168_),
    .D(_02723_),
    .X(_02814_));
 sky130_fd_sc_hd__a22o_1 _10554_ (.A1(_02993_),
    .A2(_02168_),
    .B1(_02723_),
    .B2(_00377_),
    .X(_02815_));
 sky130_fd_sc_hd__and4b_1 _10555_ (.A_N(_02814_),
    .B(_02815_),
    .C(_00095_),
    .D(_01933_),
    .X(_02816_));
 sky130_fd_sc_hd__or2_1 _10556_ (.A(_02814_),
    .B(_02816_),
    .X(_02818_));
 sky130_fd_sc_hd__and2b_1 _10557_ (.A_N(_02803_),
    .B(_02802_),
    .X(_02819_));
 sky130_fd_sc_hd__nand2_1 _10558_ (.A(_00293_),
    .B(_02169_),
    .Y(_02820_));
 sky130_fd_sc_hd__xnor2_1 _10559_ (.A(_02819_),
    .B(_02820_),
    .Y(_02821_));
 sky130_fd_sc_hd__nand2_1 _10560_ (.A(_00294_),
    .B(_01934_),
    .Y(_02822_));
 sky130_fd_sc_hd__xnor2_1 _10561_ (.A(_02818_),
    .B(_02822_),
    .Y(_02823_));
 sky130_fd_sc_hd__nand2_1 _10562_ (.A(_02821_),
    .B(_02823_),
    .Y(_02824_));
 sky130_fd_sc_hd__inv_2 _10563_ (.A(_02824_),
    .Y(_02825_));
 sky130_fd_sc_hd__a31o_1 _10564_ (.A1(_00818_),
    .A2(_02758_),
    .A3(_02818_),
    .B1(_02825_),
    .X(_02826_));
 sky130_fd_sc_hd__or2b_1 _10565_ (.A(_02804_),
    .B_N(_02801_),
    .X(_02827_));
 sky130_fd_sc_hd__nand2_1 _10566_ (.A(_02805_),
    .B(_02827_),
    .Y(_02829_));
 sky130_fd_sc_hd__xnor2_1 _10567_ (.A(_02826_),
    .B(_02829_),
    .Y(_02830_));
 sky130_fd_sc_hd__inv_2 _10568_ (.A(_02814_),
    .Y(_02831_));
 sky130_fd_sc_hd__a22oi_1 _10569_ (.A1(_00819_),
    .A2(_01934_),
    .B1(_02831_),
    .B2(_02815_),
    .Y(_02832_));
 sky130_fd_sc_hd__nor2_1 _10570_ (.A(_02816_),
    .B(_02832_),
    .Y(_02833_));
 sky130_fd_sc_hd__and4_1 _10571_ (.A(_00399_),
    .B(_03015_),
    .C(_01934_),
    .D(_02169_),
    .X(_02834_));
 sky130_fd_sc_hd__nand2_1 _10572_ (.A(_02833_),
    .B(_02834_),
    .Y(_02835_));
 sky130_fd_sc_hd__or2_1 _10573_ (.A(_02821_),
    .B(_02823_),
    .X(_02836_));
 sky130_fd_sc_hd__nand2_1 _10574_ (.A(_02824_),
    .B(_02836_),
    .Y(_02837_));
 sky130_fd_sc_hd__nor2_1 _10575_ (.A(_02835_),
    .B(_02837_),
    .Y(_02838_));
 sky130_fd_sc_hd__and2b_1 _10576_ (.A_N(_02829_),
    .B(_02826_),
    .X(_02840_));
 sky130_fd_sc_hd__a21oi_1 _10577_ (.A1(_02830_),
    .A2(_02838_),
    .B1(_02840_),
    .Y(_02841_));
 sky130_fd_sc_hd__xor2_1 _10578_ (.A(_02813_),
    .B(_02841_),
    .X(_02842_));
 sky130_fd_sc_hd__and4_1 _10579_ (.A(_00143_),
    .B(_04906_),
    .C(_02306_),
    .D(_02305_),
    .X(_02843_));
 sky130_fd_sc_hd__a22o_1 _10580_ (.A1(_00143_),
    .A2(_02306_),
    .B1(_02305_),
    .B2(_04906_),
    .X(_02844_));
 sky130_fd_sc_hd__or2b_1 _10581_ (.A(_02843_),
    .B_N(_02844_),
    .X(_02845_));
 sky130_fd_sc_hd__nand2_1 _10582_ (.A(_00310_),
    .B(_01413_),
    .Y(_02846_));
 sky130_fd_sc_hd__xnor2_1 _10583_ (.A(_02845_),
    .B(_02846_),
    .Y(_02847_));
 sky130_fd_sc_hd__a22o_1 _10584_ (.A1(_04895_),
    .A2(_02306_),
    .B1(_02305_),
    .B2(_04928_),
    .X(_02848_));
 sky130_fd_sc_hd__buf_2 _10585_ (.A(_02158_),
    .X(_02849_));
 sky130_fd_sc_hd__and4_1 _10586_ (.A(_04895_),
    .B(_04928_),
    .C(_02849_),
    .D(_02304_),
    .X(_02851_));
 sky130_fd_sc_hd__a31o_1 _10587_ (.A1(_00145_),
    .A2(_01413_),
    .A3(_02848_),
    .B1(_02851_),
    .X(_02852_));
 sky130_fd_sc_hd__or2b_1 _10588_ (.A(_02847_),
    .B_N(_02852_),
    .X(_02853_));
 sky130_fd_sc_hd__a31o_1 _10589_ (.A1(_00310_),
    .A2(_01413_),
    .A3(_02844_),
    .B1(_02843_),
    .X(_02854_));
 sky130_fd_sc_hd__clkbuf_4 _10590_ (.A(_02306_),
    .X(_02855_));
 sky130_fd_sc_hd__clkbuf_4 _10591_ (.A(_02855_),
    .X(_02856_));
 sky130_fd_sc_hd__clkbuf_4 _10592_ (.A(_02305_),
    .X(_02857_));
 sky130_fd_sc_hd__clkbuf_4 _10593_ (.A(_02857_),
    .X(_02858_));
 sky130_fd_sc_hd__nand4_1 _10594_ (.A(_00145_),
    .B(_00310_),
    .C(_02856_),
    .D(_02858_),
    .Y(_02859_));
 sky130_fd_sc_hd__a22o_1 _10595_ (.A1(_00310_),
    .A2(_02855_),
    .B1(_02857_),
    .B2(_00145_),
    .X(_02860_));
 sky130_fd_sc_hd__and3_1 _10596_ (.A(_02854_),
    .B(_02859_),
    .C(_02860_),
    .X(_02862_));
 sky130_fd_sc_hd__a21oi_1 _10597_ (.A1(_02859_),
    .A2(_02860_),
    .B1(_02854_),
    .Y(_02863_));
 sky130_fd_sc_hd__nor2_1 _10598_ (.A(_02862_),
    .B(_02863_),
    .Y(_02864_));
 sky130_fd_sc_hd__xor2_1 _10599_ (.A(_02853_),
    .B(_02864_),
    .X(_02865_));
 sky130_fd_sc_hd__and4_1 _10600_ (.A(_04862_),
    .B(_04873_),
    .C(_01410_),
    .D(_02158_),
    .X(_02866_));
 sky130_fd_sc_hd__a22o_1 _10601_ (.A1(_04862_),
    .A2(_01410_),
    .B1(_02158_),
    .B2(_04873_),
    .X(_02867_));
 sky130_fd_sc_hd__and4b_1 _10602_ (.A_N(_02866_),
    .B(_02867_),
    .C(_00142_),
    .D(_01059_),
    .X(_02868_));
 sky130_fd_sc_hd__or2_1 _10603_ (.A(_02866_),
    .B(_02868_),
    .X(_02869_));
 sky130_fd_sc_hd__and2b_1 _10604_ (.A_N(_02851_),
    .B(_02848_),
    .X(_02870_));
 sky130_fd_sc_hd__nand2_1 _10605_ (.A(_00144_),
    .B(_01412_),
    .Y(_02871_));
 sky130_fd_sc_hd__xnor2_1 _10606_ (.A(_02870_),
    .B(_02871_),
    .Y(_02873_));
 sky130_fd_sc_hd__nand2_1 _10607_ (.A(_00158_),
    .B(_01059_),
    .Y(_02874_));
 sky130_fd_sc_hd__xnor2_1 _10608_ (.A(_02869_),
    .B(_02874_),
    .Y(_02875_));
 sky130_fd_sc_hd__nand2_1 _10609_ (.A(_02873_),
    .B(_02875_),
    .Y(_02876_));
 sky130_fd_sc_hd__inv_2 _10610_ (.A(_02876_),
    .Y(_02877_));
 sky130_fd_sc_hd__a31o_1 _10611_ (.A1(_00310_),
    .A2(_01060_),
    .A3(_02869_),
    .B1(_02877_),
    .X(_02878_));
 sky130_fd_sc_hd__or2b_1 _10612_ (.A(_02852_),
    .B_N(_02847_),
    .X(_02879_));
 sky130_fd_sc_hd__nand2_1 _10613_ (.A(_02853_),
    .B(_02879_),
    .Y(_02880_));
 sky130_fd_sc_hd__or2b_1 _10614_ (.A(_02878_),
    .B_N(_02880_),
    .X(_02881_));
 sky130_fd_sc_hd__inv_2 _10615_ (.A(_02866_),
    .Y(_02882_));
 sky130_fd_sc_hd__a22oi_1 _10616_ (.A1(_01472_),
    .A2(_01060_),
    .B1(_02882_),
    .B2(_02867_),
    .Y(_02884_));
 sky130_fd_sc_hd__nor2_1 _10617_ (.A(_02868_),
    .B(_02884_),
    .Y(_02885_));
 sky130_fd_sc_hd__and4_1 _10618_ (.A(_00635_),
    .B(_04939_),
    .C(_01060_),
    .D(_01413_),
    .X(_02886_));
 sky130_fd_sc_hd__nand2_1 _10619_ (.A(_02885_),
    .B(_02886_),
    .Y(_02887_));
 sky130_fd_sc_hd__or2_1 _10620_ (.A(_02873_),
    .B(_02875_),
    .X(_02888_));
 sky130_fd_sc_hd__nand2_1 _10621_ (.A(_02876_),
    .B(_02888_),
    .Y(_02889_));
 sky130_fd_sc_hd__nor2_1 _10622_ (.A(_02887_),
    .B(_02889_),
    .Y(_02890_));
 sky130_fd_sc_hd__and2b_1 _10623_ (.A_N(_02880_),
    .B(_02878_),
    .X(_02891_));
 sky130_fd_sc_hd__a21oi_1 _10624_ (.A1(_02881_),
    .A2(_02890_),
    .B1(_02891_),
    .Y(_02892_));
 sky130_fd_sc_hd__xor2_1 _10625_ (.A(_02865_),
    .B(_02892_),
    .X(_02893_));
 sky130_fd_sc_hd__nand2_1 _10626_ (.A(_02842_),
    .B(_02893_),
    .Y(_02895_));
 sky130_fd_sc_hd__and2b_1 _10627_ (.A_N(_02805_),
    .B(_02812_),
    .X(_02896_));
 sky130_fd_sc_hd__nor2_1 _10628_ (.A(_02813_),
    .B(_02841_),
    .Y(_02897_));
 sky130_fd_sc_hd__nand2_1 _10629_ (.A(_00819_),
    .B(_02735_),
    .Y(_02898_));
 sky130_fd_sc_hd__and3_1 _10630_ (.A(_00818_),
    .B(_02731_),
    .C(_02898_),
    .X(_02899_));
 sky130_fd_sc_hd__xor2_1 _10631_ (.A(_02810_),
    .B(_02899_),
    .X(_02900_));
 sky130_fd_sc_hd__o21a_1 _10632_ (.A1(_02896_),
    .A2(_02897_),
    .B1(_02900_),
    .X(_02901_));
 sky130_fd_sc_hd__nor3_1 _10633_ (.A(_02896_),
    .B(_02897_),
    .C(_02900_),
    .Y(_02902_));
 sky130_fd_sc_hd__nor2_1 _10634_ (.A(_02901_),
    .B(_02902_),
    .Y(_02903_));
 sky130_fd_sc_hd__and2b_1 _10635_ (.A_N(_02853_),
    .B(_02864_),
    .X(_02904_));
 sky130_fd_sc_hd__nor2_1 _10636_ (.A(_02865_),
    .B(_02892_),
    .Y(_02906_));
 sky130_fd_sc_hd__nand2_1 _10637_ (.A(_01472_),
    .B(_02856_),
    .Y(_02907_));
 sky130_fd_sc_hd__and3_1 _10638_ (.A(_00859_),
    .B(_02858_),
    .C(_02907_),
    .X(_02908_));
 sky130_fd_sc_hd__xor2_1 _10639_ (.A(_02862_),
    .B(_02908_),
    .X(_02909_));
 sky130_fd_sc_hd__o21a_1 _10640_ (.A1(_02904_),
    .A2(_02906_),
    .B1(_02909_),
    .X(_02910_));
 sky130_fd_sc_hd__nor3_1 _10641_ (.A(_02904_),
    .B(_02906_),
    .C(_02909_),
    .Y(_02911_));
 sky130_fd_sc_hd__nor2_1 _10642_ (.A(_02910_),
    .B(_02911_),
    .Y(_02912_));
 sky130_fd_sc_hd__nand2_1 _10643_ (.A(_02903_),
    .B(_02912_),
    .Y(_02913_));
 sky130_fd_sc_hd__or2_1 _10644_ (.A(_02903_),
    .B(_02912_),
    .X(_02914_));
 sky130_fd_sc_hd__nand2_1 _10645_ (.A(_02913_),
    .B(_02914_),
    .Y(_02915_));
 sky130_fd_sc_hd__nor2_1 _10646_ (.A(_02895_),
    .B(_02915_),
    .Y(_02917_));
 sky130_fd_sc_hd__and2_1 _10647_ (.A(_02895_),
    .B(_02915_),
    .X(_02918_));
 sky130_fd_sc_hd__nor2_2 _10648_ (.A(_02917_),
    .B(_02918_),
    .Y(_02919_));
 sky130_fd_sc_hd__xnor2_4 _10649_ (.A(_02796_),
    .B(_02919_),
    .Y(_02920_));
 sky130_fd_sc_hd__xor2_1 _10650_ (.A(_02830_),
    .B(_02838_),
    .X(_02921_));
 sky130_fd_sc_hd__or2b_1 _10651_ (.A(_02891_),
    .B_N(_02881_),
    .X(_02922_));
 sky130_fd_sc_hd__xnor2_1 _10652_ (.A(_02922_),
    .B(_02890_),
    .Y(_02923_));
 sky130_fd_sc_hd__nand2_1 _10653_ (.A(_02921_),
    .B(_02923_),
    .Y(_02924_));
 sky130_fd_sc_hd__or2_1 _10654_ (.A(_02842_),
    .B(_02893_),
    .X(_02925_));
 sky130_fd_sc_hd__nand2_1 _10655_ (.A(_02895_),
    .B(_02925_),
    .Y(_02926_));
 sky130_fd_sc_hd__nand2_1 _10656_ (.A(_02924_),
    .B(_02926_),
    .Y(_02928_));
 sky130_fd_sc_hd__a22oi_1 _10657_ (.A1(_00636_),
    .A2(_02765_),
    .B1(_02722_),
    .B2(_01156_),
    .Y(_02929_));
 sky130_fd_sc_hd__nor2_1 _10658_ (.A(_02769_),
    .B(_02929_),
    .Y(_02930_));
 sky130_fd_sc_hd__nor2_1 _10659_ (.A(_02924_),
    .B(_02926_),
    .Y(_02931_));
 sky130_fd_sc_hd__a21o_1 _10660_ (.A1(_02928_),
    .A2(_02930_),
    .B1(_02931_),
    .X(_02932_));
 sky130_fd_sc_hd__xor2_4 _10661_ (.A(_02920_),
    .B(_02932_),
    .X(_02933_));
 sky130_fd_sc_hd__and2b_1 _10662_ (.A_N(_02931_),
    .B(_02928_),
    .X(_02934_));
 sky130_fd_sc_hd__xnor2_2 _10663_ (.A(_02930_),
    .B(_02934_),
    .Y(_02935_));
 sky130_fd_sc_hd__and2_1 _10664_ (.A(_02835_),
    .B(_02837_),
    .X(_02936_));
 sky130_fd_sc_hd__nor2_1 _10665_ (.A(_02838_),
    .B(_02936_),
    .Y(_02937_));
 sky130_fd_sc_hd__and4_1 _10666_ (.A(_00819_),
    .B(_00818_),
    .C(_02856_),
    .D(_02858_),
    .X(_02939_));
 sky130_fd_sc_hd__a22o_1 _10667_ (.A1(_05192_),
    .A2(_01546_),
    .B1(_02156_),
    .B2(_02982_),
    .X(_02940_));
 sky130_fd_sc_hd__and4_1 _10668_ (.A(_02982_),
    .B(_05192_),
    .C(_01546_),
    .D(_02156_),
    .X(_02941_));
 sky130_fd_sc_hd__a31o_1 _10669_ (.A1(_05181_),
    .A2(_01411_),
    .A3(_02940_),
    .B1(_02941_),
    .X(_02942_));
 sky130_fd_sc_hd__nand4_1 _10670_ (.A(_00094_),
    .B(_00151_),
    .C(_02849_),
    .D(_02304_),
    .Y(_02943_));
 sky130_fd_sc_hd__a22o_1 _10671_ (.A1(_05181_),
    .A2(_02849_),
    .B1(_02304_),
    .B2(_00094_),
    .X(_02944_));
 sky130_fd_sc_hd__and3_1 _10672_ (.A(_02942_),
    .B(_02943_),
    .C(_02944_),
    .X(_02945_));
 sky130_fd_sc_hd__nand2_1 _10673_ (.A(_00293_),
    .B(_02855_),
    .Y(_02946_));
 sky130_fd_sc_hd__and3_1 _10674_ (.A(_00294_),
    .B(_02857_),
    .C(_02946_),
    .X(_02947_));
 sky130_fd_sc_hd__and2_1 _10675_ (.A(_02945_),
    .B(_02947_),
    .X(_02948_));
 sky130_fd_sc_hd__or2b_1 _10676_ (.A(_02941_),
    .B_N(_02940_),
    .X(_02950_));
 sky130_fd_sc_hd__nand2_1 _10677_ (.A(_05181_),
    .B(_01411_),
    .Y(_02951_));
 sky130_fd_sc_hd__xnor2_1 _10678_ (.A(_02950_),
    .B(_02951_),
    .Y(_02952_));
 sky130_fd_sc_hd__a22o_1 _10679_ (.A1(_02982_),
    .A2(_01546_),
    .B1(_02156_),
    .B2(_00377_),
    .X(_02953_));
 sky130_fd_sc_hd__and4_1 _10680_ (.A(_00366_),
    .B(_02982_),
    .C(_01546_),
    .D(_02156_),
    .X(_02954_));
 sky130_fd_sc_hd__a31o_1 _10681_ (.A1(_00094_),
    .A2(_01411_),
    .A3(_02953_),
    .B1(_02954_),
    .X(_02955_));
 sky130_fd_sc_hd__and2b_1 _10682_ (.A_N(_02952_),
    .B(_02955_),
    .X(_02956_));
 sky130_fd_sc_hd__a21oi_1 _10683_ (.A1(_02943_),
    .A2(_02944_),
    .B1(_02942_),
    .Y(_02957_));
 sky130_fd_sc_hd__nor2_1 _10684_ (.A(_02945_),
    .B(_02957_),
    .Y(_02958_));
 sky130_fd_sc_hd__and2_1 _10685_ (.A(_02956_),
    .B(_02958_),
    .X(_02959_));
 sky130_fd_sc_hd__nand2_1 _10686_ (.A(_05181_),
    .B(_01058_),
    .Y(_02961_));
 sky130_fd_sc_hd__a22o_1 _10687_ (.A1(_02982_),
    .A2(net50),
    .B1(_02158_),
    .B2(_00366_),
    .X(_02962_));
 sky130_fd_sc_hd__and4_1 _10688_ (.A(_00366_),
    .B(_02982_),
    .C(net50),
    .D(_01546_),
    .X(_02963_));
 sky130_fd_sc_hd__a31o_1 _10689_ (.A1(_05203_),
    .A2(_01058_),
    .A3(_02962_),
    .B1(_02963_),
    .X(_02964_));
 sky130_fd_sc_hd__or2b_1 _10690_ (.A(_02961_),
    .B_N(_02964_),
    .X(_02965_));
 sky130_fd_sc_hd__and2b_1 _10691_ (.A_N(_02954_),
    .B(_02953_),
    .X(_02966_));
 sky130_fd_sc_hd__nand2_1 _10692_ (.A(_00094_),
    .B(_01411_),
    .Y(_02967_));
 sky130_fd_sc_hd__xnor2_1 _10693_ (.A(_02966_),
    .B(_02967_),
    .Y(_02968_));
 sky130_fd_sc_hd__xnor2_1 _10694_ (.A(_02964_),
    .B(_02961_),
    .Y(_02969_));
 sky130_fd_sc_hd__nand2_1 _10695_ (.A(_02968_),
    .B(_02969_),
    .Y(_02970_));
 sky130_fd_sc_hd__xor2_1 _10696_ (.A(_02955_),
    .B(_02952_),
    .X(_02972_));
 sky130_fd_sc_hd__a21o_1 _10697_ (.A1(_02965_),
    .A2(_02970_),
    .B1(_02972_),
    .X(_02973_));
 sky130_fd_sc_hd__nand3_1 _10698_ (.A(_02965_),
    .B(_02970_),
    .C(_02972_),
    .Y(_02974_));
 sky130_fd_sc_hd__nand2_1 _10699_ (.A(_02973_),
    .B(_02974_),
    .Y(_02975_));
 sky130_fd_sc_hd__and2b_1 _10700_ (.A_N(_02963_),
    .B(_02962_),
    .X(_02976_));
 sky130_fd_sc_hd__nand2_1 _10701_ (.A(_00095_),
    .B(_01059_),
    .Y(_02977_));
 sky130_fd_sc_hd__xnor2_1 _10702_ (.A(_02976_),
    .B(_02977_),
    .Y(_02978_));
 sky130_fd_sc_hd__and4_1 _10703_ (.A(_00388_),
    .B(_03004_),
    .C(_01059_),
    .D(_01412_),
    .X(_02979_));
 sky130_fd_sc_hd__nand2_1 _10704_ (.A(_02978_),
    .B(_02979_),
    .Y(_02980_));
 sky130_fd_sc_hd__or2_1 _10705_ (.A(_02968_),
    .B(_02969_),
    .X(_02981_));
 sky130_fd_sc_hd__nand2_1 _10706_ (.A(_02970_),
    .B(_02981_),
    .Y(_02983_));
 sky130_fd_sc_hd__or3_1 _10707_ (.A(_02975_),
    .B(_02980_),
    .C(_02983_),
    .X(_02984_));
 sky130_fd_sc_hd__nor2_1 _10708_ (.A(_02956_),
    .B(_02958_),
    .Y(_02985_));
 sky130_fd_sc_hd__or2_1 _10709_ (.A(_02959_),
    .B(_02985_),
    .X(_02986_));
 sky130_fd_sc_hd__a21oi_1 _10710_ (.A1(_02973_),
    .A2(_02984_),
    .B1(_02986_),
    .Y(_02987_));
 sky130_fd_sc_hd__xor2_1 _10711_ (.A(_02945_),
    .B(_02947_),
    .X(_02988_));
 sky130_fd_sc_hd__o21a_1 _10712_ (.A1(_02959_),
    .A2(_02987_),
    .B1(_02988_),
    .X(_02989_));
 sky130_fd_sc_hd__or4_1 _10713_ (.A(_02937_),
    .B(_02939_),
    .C(_02948_),
    .D(_02989_),
    .X(_02990_));
 sky130_fd_sc_hd__o31ai_2 _10714_ (.A1(_02939_),
    .A2(_02948_),
    .A3(_02989_),
    .B1(_02937_),
    .Y(_02991_));
 sky130_fd_sc_hd__and2_1 _10715_ (.A(_02887_),
    .B(_02889_),
    .X(_02992_));
 sky130_fd_sc_hd__or2_1 _10716_ (.A(_02890_),
    .B(_02992_),
    .X(_02994_));
 sky130_fd_sc_hd__nand2_1 _10717_ (.A(_02991_),
    .B(_02994_),
    .Y(_02995_));
 sky130_fd_sc_hd__or2_1 _10718_ (.A(_02921_),
    .B(_02923_),
    .X(_02996_));
 sky130_fd_sc_hd__and2_1 _10719_ (.A(_02924_),
    .B(_02996_),
    .X(_02997_));
 sky130_fd_sc_hd__a21oi_1 _10720_ (.A1(_02990_),
    .A2(_02995_),
    .B1(_02997_),
    .Y(_02998_));
 sky130_fd_sc_hd__and3_1 _10721_ (.A(_02997_),
    .B(_02990_),
    .C(_02995_),
    .X(_02999_));
 sky130_fd_sc_hd__a21oi_1 _10722_ (.A1(_01156_),
    .A2(_02766_),
    .B1(_02999_),
    .Y(_03000_));
 sky130_fd_sc_hd__or2_2 _10723_ (.A(_02998_),
    .B(_03000_),
    .X(_03001_));
 sky130_fd_sc_hd__xor2_1 _10724_ (.A(_02935_),
    .B(_03001_),
    .X(_03002_));
 sky130_fd_sc_hd__inv_2 _10725_ (.A(_03002_),
    .Y(_03003_));
 sky130_fd_sc_hd__nand2_1 _10726_ (.A(_02990_),
    .B(_02991_),
    .Y(_03005_));
 sky130_fd_sc_hd__xor2_1 _10727_ (.A(_02994_),
    .B(_03005_),
    .X(_03006_));
 sky130_fd_sc_hd__or2_1 _10728_ (.A(_02833_),
    .B(_02834_),
    .X(_03007_));
 sky130_fd_sc_hd__nand2_1 _10729_ (.A(_02835_),
    .B(_03007_),
    .Y(_03008_));
 sky130_fd_sc_hd__nor3_1 _10730_ (.A(_02988_),
    .B(_02959_),
    .C(_02987_),
    .Y(_03009_));
 sky130_fd_sc_hd__or2_1 _10731_ (.A(_02989_),
    .B(_03009_),
    .X(_03010_));
 sky130_fd_sc_hd__nand2_1 _10732_ (.A(_03008_),
    .B(_03010_),
    .Y(_03011_));
 sky130_fd_sc_hd__or2_1 _10733_ (.A(_02885_),
    .B(_02886_),
    .X(_03012_));
 sky130_fd_sc_hd__nand2_1 _10734_ (.A(_02887_),
    .B(_03012_),
    .Y(_03013_));
 sky130_fd_sc_hd__o21ai_1 _10735_ (.A1(_03008_),
    .A2(_03010_),
    .B1(_03013_),
    .Y(_03014_));
 sky130_fd_sc_hd__and3_1 _10736_ (.A(_03006_),
    .B(_03011_),
    .C(_03014_),
    .X(_03016_));
 sky130_fd_sc_hd__nand4_1 _10737_ (.A(_00399_),
    .B(_03015_),
    .C(_02758_),
    .D(_02721_),
    .Y(_03017_));
 sky130_fd_sc_hd__a22o_1 _10738_ (.A1(_03015_),
    .A2(_02758_),
    .B1(_02720_),
    .B2(_00399_),
    .X(_03018_));
 sky130_fd_sc_hd__and3_1 _10739_ (.A(_02986_),
    .B(_02973_),
    .C(_02984_),
    .X(_03019_));
 sky130_fd_sc_hd__nor2_1 _10740_ (.A(_02987_),
    .B(_03019_),
    .Y(_03020_));
 sky130_fd_sc_hd__a21oi_1 _10741_ (.A1(_03017_),
    .A2(_03018_),
    .B1(_03020_),
    .Y(_03021_));
 sky130_fd_sc_hd__a22oi_1 _10742_ (.A1(_00635_),
    .A2(_01061_),
    .B1(_01414_),
    .B2(_07040_),
    .Y(_03022_));
 sky130_fd_sc_hd__or2_1 _10743_ (.A(_02886_),
    .B(_03022_),
    .X(_03023_));
 sky130_fd_sc_hd__and3_1 _10744_ (.A(_03017_),
    .B(_03018_),
    .C(_03020_),
    .X(_03024_));
 sky130_fd_sc_hd__o21bai_1 _10745_ (.A1(_03021_),
    .A2(_03023_),
    .B1_N(_03024_),
    .Y(_03025_));
 sky130_fd_sc_hd__xor2_1 _10746_ (.A(_03008_),
    .B(_03010_),
    .X(_03027_));
 sky130_fd_sc_hd__xnor2_1 _10747_ (.A(_03013_),
    .B(_03027_),
    .Y(_03028_));
 sky130_fd_sc_hd__and2_1 _10748_ (.A(_03025_),
    .B(_03028_),
    .X(_03029_));
 sky130_fd_sc_hd__nor2_1 _10749_ (.A(_03025_),
    .B(_03028_),
    .Y(_03030_));
 sky130_fd_sc_hd__or2_1 _10750_ (.A(_03029_),
    .B(_03030_),
    .X(_03031_));
 sky130_fd_sc_hd__nor2_1 _10751_ (.A(_02980_),
    .B(_02983_),
    .Y(_03032_));
 sky130_fd_sc_hd__xnor2_1 _10752_ (.A(_02975_),
    .B(_03032_),
    .Y(_03033_));
 sky130_fd_sc_hd__a21o_1 _10753_ (.A1(_00399_),
    .A2(_02765_),
    .B1(_03033_),
    .X(_03034_));
 sky130_fd_sc_hd__and3_1 _10754_ (.A(_00399_),
    .B(_02759_),
    .C(_03033_),
    .X(_03035_));
 sky130_fd_sc_hd__a21o_1 _10755_ (.A1(_00526_),
    .A2(_01061_),
    .B1(_03035_),
    .X(_03036_));
 sky130_fd_sc_hd__nand2_1 _10756_ (.A(_03034_),
    .B(_03036_),
    .Y(_03038_));
 sky130_fd_sc_hd__or2_1 _10757_ (.A(_03024_),
    .B(_03021_),
    .X(_03039_));
 sky130_fd_sc_hd__xnor2_1 _10758_ (.A(_03023_),
    .B(_03039_),
    .Y(_03040_));
 sky130_fd_sc_hd__nor2_1 _10759_ (.A(_03038_),
    .B(_03040_),
    .Y(_03041_));
 sky130_fd_sc_hd__and2b_1 _10760_ (.A_N(_03031_),
    .B(_03041_),
    .X(_03042_));
 sky130_fd_sc_hd__a21oi_1 _10761_ (.A1(_03011_),
    .A2(_03014_),
    .B1(_03006_),
    .Y(_03043_));
 sky130_fd_sc_hd__nor2_1 _10762_ (.A(_03016_),
    .B(_03043_),
    .Y(_03044_));
 sky130_fd_sc_hd__o21a_1 _10763_ (.A1(_03029_),
    .A2(_03042_),
    .B1(_03044_),
    .X(_03045_));
 sky130_fd_sc_hd__o211ai_1 _10764_ (.A1(_02998_),
    .A2(_02999_),
    .B1(_01156_),
    .C1(_02766_),
    .Y(_03046_));
 sky130_fd_sc_hd__a211o_1 _10765_ (.A1(_01156_),
    .A2(_02766_),
    .B1(_02998_),
    .C1(_02999_),
    .X(_03047_));
 sky130_fd_sc_hd__nand2_1 _10766_ (.A(_03046_),
    .B(_03047_),
    .Y(_03049_));
 sky130_fd_sc_hd__o21ai_1 _10767_ (.A1(_03016_),
    .A2(_03045_),
    .B1(_03049_),
    .Y(_03050_));
 sky130_fd_sc_hd__nor2_1 _10768_ (.A(_03003_),
    .B(_03050_),
    .Y(_03051_));
 sky130_fd_sc_hd__o21bai_4 _10769_ (.A1(_02935_),
    .A2(_03001_),
    .B1_N(_03051_),
    .Y(_03052_));
 sky130_fd_sc_hd__xnor2_4 _10770_ (.A(_02933_),
    .B(_03052_),
    .Y(_03053_));
 sky130_fd_sc_hd__and4_1 _10771_ (.A(_02160_),
    .B(_06461_),
    .C(_02724_),
    .D(_02727_),
    .X(_03054_));
 sky130_fd_sc_hd__a22o_1 _10772_ (.A1(_06461_),
    .A2(_02724_),
    .B1(_02727_),
    .B2(_02160_),
    .X(_03055_));
 sky130_fd_sc_hd__or2b_1 _10773_ (.A(_03054_),
    .B_N(_03055_),
    .X(_03056_));
 sky130_fd_sc_hd__nand2_1 _10774_ (.A(_06494_),
    .B(_02168_),
    .Y(_03057_));
 sky130_fd_sc_hd__xnor2_1 _10775_ (.A(_03056_),
    .B(_03057_),
    .Y(_03058_));
 sky130_fd_sc_hd__a22o_1 _10776_ (.A1(_02160_),
    .A2(_02723_),
    .B1(_02727_),
    .B2(_02116_),
    .X(_03060_));
 sky130_fd_sc_hd__and4_1 _10777_ (.A(_02116_),
    .B(_02149_),
    .C(_02723_),
    .D(_02727_),
    .X(_03061_));
 sky130_fd_sc_hd__a31o_1 _10778_ (.A1(_06937_),
    .A2(_02169_),
    .A3(_03060_),
    .B1(_03061_),
    .X(_03062_));
 sky130_fd_sc_hd__or2b_1 _10779_ (.A(_03058_),
    .B_N(_03062_),
    .X(_03063_));
 sky130_fd_sc_hd__a31o_1 _10780_ (.A1(_06637_),
    .A2(_02720_),
    .A3(_03055_),
    .B1(_03054_),
    .X(_03064_));
 sky130_fd_sc_hd__and4_1 _10781_ (.A(_06937_),
    .B(_06494_),
    .C(_02725_),
    .D(_02730_),
    .X(_03065_));
 sky130_fd_sc_hd__a22oi_1 _10782_ (.A1(_06637_),
    .A2(_02726_),
    .B1(_02730_),
    .B2(_06937_),
    .Y(_03066_));
 sky130_fd_sc_hd__nor2_1 _10783_ (.A(_03065_),
    .B(_03066_),
    .Y(_03067_));
 sky130_fd_sc_hd__nand2_1 _10784_ (.A(_03064_),
    .B(_03067_),
    .Y(_03068_));
 sky130_fd_sc_hd__or2_1 _10785_ (.A(_03064_),
    .B(_03067_),
    .X(_03069_));
 sky130_fd_sc_hd__and2_1 _10786_ (.A(_03068_),
    .B(_03069_),
    .X(_03071_));
 sky130_fd_sc_hd__and2b_1 _10787_ (.A_N(_03063_),
    .B(_03071_),
    .X(_03072_));
 sky130_fd_sc_hd__xor2_1 _10788_ (.A(_03063_),
    .B(_03071_),
    .X(_03073_));
 sky130_fd_sc_hd__and4_1 _10789_ (.A(_00628_),
    .B(_00650_),
    .C(net54),
    .D(_02312_),
    .X(_03074_));
 sky130_fd_sc_hd__inv_2 _10790_ (.A(_03074_),
    .Y(_03075_));
 sky130_fd_sc_hd__a22o_1 _10791_ (.A1(_02149_),
    .A2(net54),
    .B1(_02312_),
    .B2(_02105_),
    .X(_03076_));
 sky130_fd_sc_hd__and4_1 _10792_ (.A(_05588_),
    .B(_01933_),
    .C(_03075_),
    .D(_03076_),
    .X(_03077_));
 sky130_fd_sc_hd__a22oi_1 _10793_ (.A1(_06937_),
    .A2(_02758_),
    .B1(_03075_),
    .B2(_03076_),
    .Y(_03078_));
 sky130_fd_sc_hd__nor2_1 _10794_ (.A(_03077_),
    .B(_03078_),
    .Y(_03079_));
 sky130_fd_sc_hd__and4_1 _10795_ (.A(_02259_),
    .B(_02171_),
    .C(_02758_),
    .D(_02169_),
    .X(_03080_));
 sky130_fd_sc_hd__nand2_1 _10796_ (.A(_03079_),
    .B(_03080_),
    .Y(_03082_));
 sky130_fd_sc_hd__and2b_1 _10797_ (.A_N(_03061_),
    .B(_03060_),
    .X(_03083_));
 sky130_fd_sc_hd__nand2_1 _10798_ (.A(_06461_),
    .B(_02168_),
    .Y(_03084_));
 sky130_fd_sc_hd__xnor2_1 _10799_ (.A(_03083_),
    .B(_03084_),
    .Y(_03085_));
 sky130_fd_sc_hd__or2_1 _10800_ (.A(_03074_),
    .B(_03077_),
    .X(_03086_));
 sky130_fd_sc_hd__nand2_1 _10801_ (.A(_06483_),
    .B(_01933_),
    .Y(_03087_));
 sky130_fd_sc_hd__xnor2_1 _10802_ (.A(_03086_),
    .B(_03087_),
    .Y(_03088_));
 sky130_fd_sc_hd__nand2_1 _10803_ (.A(_03085_),
    .B(_03088_),
    .Y(_03089_));
 sky130_fd_sc_hd__or2_1 _10804_ (.A(_03085_),
    .B(_03088_),
    .X(_03090_));
 sky130_fd_sc_hd__nand2_1 _10805_ (.A(_03089_),
    .B(_03090_),
    .Y(_03091_));
 sky130_fd_sc_hd__nor2_1 _10806_ (.A(_03082_),
    .B(_03091_),
    .Y(_03093_));
 sky130_fd_sc_hd__inv_2 _10807_ (.A(_03089_),
    .Y(_03094_));
 sky130_fd_sc_hd__a31o_1 _10808_ (.A1(_06494_),
    .A2(_01934_),
    .A3(_03086_),
    .B1(_03094_),
    .X(_03095_));
 sky130_fd_sc_hd__or2b_1 _10809_ (.A(_03062_),
    .B_N(_03058_),
    .X(_03096_));
 sky130_fd_sc_hd__nand2_1 _10810_ (.A(_03063_),
    .B(_03096_),
    .Y(_03097_));
 sky130_fd_sc_hd__or2b_1 _10811_ (.A(_03095_),
    .B_N(_03097_),
    .X(_03098_));
 sky130_fd_sc_hd__and2b_1 _10812_ (.A_N(_03097_),
    .B(_03095_),
    .X(_03099_));
 sky130_fd_sc_hd__a21oi_1 _10813_ (.A1(_03093_),
    .A2(_03098_),
    .B1(_03099_),
    .Y(_03100_));
 sky130_fd_sc_hd__nor2_1 _10814_ (.A(_03073_),
    .B(_03100_),
    .Y(_03101_));
 sky130_fd_sc_hd__nand2_1 _10815_ (.A(_06937_),
    .B(_02735_),
    .Y(_03102_));
 sky130_fd_sc_hd__and3_1 _10816_ (.A(_06637_),
    .B(_02731_),
    .C(_03102_),
    .X(_03104_));
 sky130_fd_sc_hd__xnor2_1 _10817_ (.A(_03068_),
    .B(_03104_),
    .Y(_03105_));
 sky130_fd_sc_hd__o21a_1 _10818_ (.A1(_03072_),
    .A2(_03101_),
    .B1(_03105_),
    .X(_03106_));
 sky130_fd_sc_hd__nor3_1 _10819_ (.A(_03105_),
    .B(_03072_),
    .C(_03101_),
    .Y(_03107_));
 sky130_fd_sc_hd__nor2_1 _10820_ (.A(_03106_),
    .B(_03107_),
    .Y(_03108_));
 sky130_fd_sc_hd__a22o_1 _10821_ (.A1(_00891_),
    .A2(net56),
    .B1(net57),
    .B2(_00989_),
    .X(_03109_));
 sky130_fd_sc_hd__and4_1 _10822_ (.A(_03587_),
    .B(_00891_),
    .C(net56),
    .D(net57),
    .X(_03110_));
 sky130_fd_sc_hd__a31oi_2 _10823_ (.A1(_01339_),
    .A2(net54),
    .A3(_03109_),
    .B1(_03110_),
    .Y(_03111_));
 sky130_fd_sc_hd__and4_1 _10824_ (.A(_01372_),
    .B(_04268_),
    .C(_02312_),
    .D(net57),
    .X(_03112_));
 sky130_fd_sc_hd__a22oi_1 _10825_ (.A1(_01339_),
    .A2(_02312_),
    .B1(net57),
    .B2(_04081_),
    .Y(_03113_));
 sky130_fd_sc_hd__or2_1 _10826_ (.A(_03112_),
    .B(_03113_),
    .X(_03115_));
 sky130_fd_sc_hd__nor2_1 _10827_ (.A(_03111_),
    .B(_03115_),
    .Y(_03116_));
 sky130_fd_sc_hd__nand2_1 _10828_ (.A(_01383_),
    .B(_02724_),
    .Y(_03117_));
 sky130_fd_sc_hd__and3_1 _10829_ (.A(_01350_),
    .B(_02728_),
    .C(_03117_),
    .X(_03118_));
 sky130_fd_sc_hd__a32o_1 _10830_ (.A1(_04081_),
    .A2(net54),
    .A3(_02508_),
    .B1(_02507_),
    .B2(_02727_),
    .X(_03119_));
 sky130_fd_sc_hd__and2b_1 _10831_ (.A_N(_03110_),
    .B(_03109_),
    .X(_03120_));
 sky130_fd_sc_hd__nand2_1 _10832_ (.A(_01339_),
    .B(net54),
    .Y(_03121_));
 sky130_fd_sc_hd__xnor2_2 _10833_ (.A(_03120_),
    .B(_03121_),
    .Y(_03122_));
 sky130_fd_sc_hd__xor2_1 _10834_ (.A(_03111_),
    .B(_03115_),
    .X(_03123_));
 sky130_fd_sc_hd__and3_1 _10835_ (.A(_03119_),
    .B(_03122_),
    .C(_03123_),
    .X(_03124_));
 sky130_fd_sc_hd__and3_1 _10836_ (.A(_01339_),
    .B(_01933_),
    .C(_02513_),
    .X(_03126_));
 sky130_fd_sc_hd__a21o_1 _10837_ (.A1(_02512_),
    .A2(_02515_),
    .B1(_03126_),
    .X(_03127_));
 sky130_fd_sc_hd__xor2_1 _10838_ (.A(_03119_),
    .B(_03122_),
    .X(_03128_));
 sky130_fd_sc_hd__and2_1 _10839_ (.A(_03127_),
    .B(_03128_),
    .X(_03129_));
 sky130_fd_sc_hd__xnor2_1 _10840_ (.A(_03127_),
    .B(_03128_),
    .Y(_03130_));
 sky130_fd_sc_hd__nor2_1 _10841_ (.A(_02517_),
    .B(_03130_),
    .Y(_03131_));
 sky130_fd_sc_hd__a21oi_1 _10842_ (.A1(_03119_),
    .A2(_03122_),
    .B1(_03123_),
    .Y(_03132_));
 sky130_fd_sc_hd__nor2_1 _10843_ (.A(_03124_),
    .B(_03132_),
    .Y(_03133_));
 sky130_fd_sc_hd__o21a_1 _10844_ (.A1(_03129_),
    .A2(_03131_),
    .B1(_03133_),
    .X(_03134_));
 sky130_fd_sc_hd__xor2_1 _10845_ (.A(_03116_),
    .B(_03118_),
    .X(_03135_));
 sky130_fd_sc_hd__o21a_1 _10846_ (.A1(_03124_),
    .A2(_03134_),
    .B1(_03135_),
    .X(_03137_));
 sky130_fd_sc_hd__a211o_1 _10847_ (.A1(_03116_),
    .A2(_03118_),
    .B1(_03137_),
    .C1(_03112_),
    .X(_03138_));
 sky130_fd_sc_hd__a22o_1 _10848_ (.A1(_00541_),
    .A2(_01545_),
    .B1(net52),
    .B2(_05742_),
    .X(_03139_));
 sky130_fd_sc_hd__and4_1 _10849_ (.A(_05742_),
    .B(_00541_),
    .C(_01545_),
    .D(net52),
    .X(_03140_));
 sky130_fd_sc_hd__a31oi_2 _10850_ (.A1(_05566_),
    .A2(_01410_),
    .A3(_03139_),
    .B1(_03140_),
    .Y(_03141_));
 sky130_fd_sc_hd__and4_1 _10851_ (.A(_02664_),
    .B(_03268_),
    .C(_01546_),
    .D(_02156_),
    .X(_03142_));
 sky130_fd_sc_hd__a22oi_1 _10852_ (.A1(_03268_),
    .A2(_02158_),
    .B1(_02304_),
    .B2(_05577_),
    .Y(_03143_));
 sky130_fd_sc_hd__or2_1 _10853_ (.A(_03142_),
    .B(_03143_),
    .X(_03144_));
 sky130_fd_sc_hd__nor2_1 _10854_ (.A(_03141_),
    .B(_03144_),
    .Y(_03145_));
 sky130_fd_sc_hd__nand2_1 _10855_ (.A(_06461_),
    .B(_02855_),
    .Y(_03146_));
 sky130_fd_sc_hd__and3_1 _10856_ (.A(_06483_),
    .B(_02857_),
    .C(_03146_),
    .X(_03148_));
 sky130_fd_sc_hd__a32o_1 _10857_ (.A1(_05588_),
    .A2(_01410_),
    .A3(_02525_),
    .B1(_02524_),
    .B2(_02304_),
    .X(_03149_));
 sky130_fd_sc_hd__and2b_1 _10858_ (.A_N(_03140_),
    .B(_03139_),
    .X(_03150_));
 sky130_fd_sc_hd__nand2_1 _10859_ (.A(_03268_),
    .B(_01410_),
    .Y(_03151_));
 sky130_fd_sc_hd__xnor2_2 _10860_ (.A(_03150_),
    .B(_03151_),
    .Y(_03152_));
 sky130_fd_sc_hd__xor2_1 _10861_ (.A(_03141_),
    .B(_03144_),
    .X(_03153_));
 sky130_fd_sc_hd__and3_1 _10862_ (.A(_03149_),
    .B(_03152_),
    .C(_03153_),
    .X(_03154_));
 sky130_fd_sc_hd__and3_1 _10863_ (.A(_05566_),
    .B(_01058_),
    .C(_02529_),
    .X(_03155_));
 sky130_fd_sc_hd__a21o_1 _10864_ (.A1(_02528_),
    .A2(_02531_),
    .B1(_03155_),
    .X(_03156_));
 sky130_fd_sc_hd__xor2_1 _10865_ (.A(_03149_),
    .B(_03152_),
    .X(_03157_));
 sky130_fd_sc_hd__and2_1 _10866_ (.A(_03156_),
    .B(_03157_),
    .X(_03159_));
 sky130_fd_sc_hd__xnor2_1 _10867_ (.A(_03156_),
    .B(_03157_),
    .Y(_03160_));
 sky130_fd_sc_hd__nor2_1 _10868_ (.A(_02534_),
    .B(_03160_),
    .Y(_03161_));
 sky130_fd_sc_hd__a21oi_1 _10869_ (.A1(_03149_),
    .A2(_03152_),
    .B1(_03153_),
    .Y(_03162_));
 sky130_fd_sc_hd__nor2_1 _10870_ (.A(_03154_),
    .B(_03162_),
    .Y(_03163_));
 sky130_fd_sc_hd__o21a_1 _10871_ (.A1(_03159_),
    .A2(_03161_),
    .B1(_03163_),
    .X(_03164_));
 sky130_fd_sc_hd__xor2_1 _10872_ (.A(_03145_),
    .B(_03148_),
    .X(_03165_));
 sky130_fd_sc_hd__o21a_1 _10873_ (.A1(_03154_),
    .A2(_03164_),
    .B1(_03165_),
    .X(_03166_));
 sky130_fd_sc_hd__a211o_1 _10874_ (.A1(_03145_),
    .A2(_03148_),
    .B1(_03166_),
    .C1(_03142_),
    .X(_03167_));
 sky130_fd_sc_hd__and2_1 _10875_ (.A(_03138_),
    .B(_03167_),
    .X(_03168_));
 sky130_fd_sc_hd__or2b_1 _10876_ (.A(_03099_),
    .B_N(_03098_),
    .X(_03170_));
 sky130_fd_sc_hd__xnor2_1 _10877_ (.A(_03093_),
    .B(_03170_),
    .Y(_03171_));
 sky130_fd_sc_hd__and2_1 _10878_ (.A(_03168_),
    .B(_03171_),
    .X(_03172_));
 sky130_fd_sc_hd__nor2_1 _10879_ (.A(_03168_),
    .B(_03171_),
    .Y(_03173_));
 sky130_fd_sc_hd__or2_1 _10880_ (.A(_03172_),
    .B(_03173_),
    .X(_03174_));
 sky130_fd_sc_hd__and2_1 _10881_ (.A(_03082_),
    .B(_03091_),
    .X(_03175_));
 sky130_fd_sc_hd__nor2_1 _10882_ (.A(_03093_),
    .B(_03175_),
    .Y(_03176_));
 sky130_fd_sc_hd__nor3_1 _10883_ (.A(_03135_),
    .B(_03124_),
    .C(_03134_),
    .Y(_03177_));
 sky130_fd_sc_hd__nor2_1 _10884_ (.A(_03137_),
    .B(_03177_),
    .Y(_03178_));
 sky130_fd_sc_hd__nor3_1 _10885_ (.A(_03165_),
    .B(_03154_),
    .C(_03164_),
    .Y(_03179_));
 sky130_fd_sc_hd__nor2_1 _10886_ (.A(_03166_),
    .B(_03179_),
    .Y(_03181_));
 sky130_fd_sc_hd__nand2_1 _10887_ (.A(_03178_),
    .B(_03181_),
    .Y(_03182_));
 sky130_fd_sc_hd__xnor2_1 _10888_ (.A(_03138_),
    .B(_03167_),
    .Y(_03183_));
 sky130_fd_sc_hd__nand2_1 _10889_ (.A(_03182_),
    .B(_03183_),
    .Y(_03184_));
 sky130_fd_sc_hd__nor2_1 _10890_ (.A(_03182_),
    .B(_03183_),
    .Y(_03185_));
 sky130_fd_sc_hd__a21oi_1 _10891_ (.A1(_03176_),
    .A2(_03184_),
    .B1(_03185_),
    .Y(_03186_));
 sky130_fd_sc_hd__nor2_1 _10892_ (.A(_03174_),
    .B(_03186_),
    .Y(_03187_));
 sky130_fd_sc_hd__and2_1 _10893_ (.A(_03174_),
    .B(_03186_),
    .X(_03188_));
 sky130_fd_sc_hd__nor2_1 _10894_ (.A(_03187_),
    .B(_03188_),
    .Y(_03189_));
 sky130_fd_sc_hd__and2b_1 _10895_ (.A_N(_03185_),
    .B(_03184_),
    .X(_03190_));
 sky130_fd_sc_hd__xor2_1 _10896_ (.A(_03176_),
    .B(_03190_),
    .X(_03192_));
 sky130_fd_sc_hd__nor3_1 _10897_ (.A(_03133_),
    .B(_03129_),
    .C(_03131_),
    .Y(_03193_));
 sky130_fd_sc_hd__nor2_1 _10898_ (.A(_03134_),
    .B(_03193_),
    .Y(_03194_));
 sky130_fd_sc_hd__nor3_1 _10899_ (.A(_03163_),
    .B(_03159_),
    .C(_03161_),
    .Y(_03195_));
 sky130_fd_sc_hd__nor2_1 _10900_ (.A(_03164_),
    .B(_03195_),
    .Y(_03196_));
 sky130_fd_sc_hd__nand2_1 _10901_ (.A(_03194_),
    .B(_03196_),
    .Y(_03197_));
 sky130_fd_sc_hd__xnor2_1 _10902_ (.A(_03178_),
    .B(_03181_),
    .Y(_03198_));
 sky130_fd_sc_hd__nor2_1 _10903_ (.A(_03197_),
    .B(_03198_),
    .Y(_03199_));
 sky130_fd_sc_hd__or2_1 _10904_ (.A(_03079_),
    .B(_03080_),
    .X(_03200_));
 sky130_fd_sc_hd__nand2_1 _10905_ (.A(_03082_),
    .B(_03200_),
    .Y(_03201_));
 sky130_fd_sc_hd__and2_1 _10906_ (.A(_03197_),
    .B(_03198_),
    .X(_03203_));
 sky130_fd_sc_hd__nor2_1 _10907_ (.A(_03201_),
    .B(_03203_),
    .Y(_03204_));
 sky130_fd_sc_hd__or3_2 _10908_ (.A(_03192_),
    .B(_03199_),
    .C(_03204_),
    .X(_03205_));
 sky130_fd_sc_hd__nor2_1 _10909_ (.A(_03199_),
    .B(_03203_),
    .Y(_03206_));
 sky130_fd_sc_hd__xnor2_2 _10910_ (.A(_03201_),
    .B(_03206_),
    .Y(_03207_));
 sky130_fd_sc_hd__and2_1 _10911_ (.A(_02517_),
    .B(_03130_),
    .X(_03208_));
 sky130_fd_sc_hd__nor2_1 _10912_ (.A(_03131_),
    .B(_03208_),
    .Y(_03209_));
 sky130_fd_sc_hd__and2_1 _10913_ (.A(_02534_),
    .B(_03160_),
    .X(_03210_));
 sky130_fd_sc_hd__nor2_1 _10914_ (.A(_03161_),
    .B(_03210_),
    .Y(_03211_));
 sky130_fd_sc_hd__nand2_1 _10915_ (.A(_03209_),
    .B(_03211_),
    .Y(_03212_));
 sky130_fd_sc_hd__xnor2_1 _10916_ (.A(_03194_),
    .B(_03196_),
    .Y(_03214_));
 sky130_fd_sc_hd__nor2_1 _10917_ (.A(_03212_),
    .B(_03214_),
    .Y(_03215_));
 sky130_fd_sc_hd__and2_1 _10918_ (.A(_03212_),
    .B(_03214_),
    .X(_03216_));
 sky130_fd_sc_hd__a22oi_1 _10919_ (.A1(_02171_),
    .A2(_02758_),
    .B1(_02720_),
    .B2(_02467_),
    .Y(_03217_));
 sky130_fd_sc_hd__nor2_1 _10920_ (.A(_03080_),
    .B(_03217_),
    .Y(_03218_));
 sky130_fd_sc_hd__and2b_1 _10921_ (.A_N(_03216_),
    .B(_03218_),
    .X(_03219_));
 sky130_fd_sc_hd__nor2_1 _10922_ (.A(_03215_),
    .B(_03219_),
    .Y(_03220_));
 sky130_fd_sc_hd__xnor2_2 _10923_ (.A(_03207_),
    .B(_03220_),
    .Y(_03221_));
 sky130_fd_sc_hd__or2_1 _10924_ (.A(_03215_),
    .B(_03216_),
    .X(_03222_));
 sky130_fd_sc_hd__xnor2_1 _10925_ (.A(_03218_),
    .B(_03222_),
    .Y(_03223_));
 sky130_fd_sc_hd__and2_1 _10926_ (.A(_02467_),
    .B(_02758_),
    .X(_03225_));
 sky130_fd_sc_hd__and2_1 _10927_ (.A(_02522_),
    .B(_02536_),
    .X(_03226_));
 sky130_fd_sc_hd__or2_1 _10928_ (.A(_03209_),
    .B(_03211_),
    .X(_03227_));
 sky130_fd_sc_hd__nand2_1 _10929_ (.A(_03212_),
    .B(_03227_),
    .Y(_03228_));
 sky130_fd_sc_hd__nor3_1 _10930_ (.A(_02520_),
    .B(_03226_),
    .C(_03228_),
    .Y(_03229_));
 sky130_fd_sc_hd__o21a_1 _10931_ (.A1(_02520_),
    .A2(_03226_),
    .B1(_03228_),
    .X(_03230_));
 sky130_fd_sc_hd__o21bai_1 _10932_ (.A1(_03225_),
    .A2(_03229_),
    .B1_N(_03230_),
    .Y(_03231_));
 sky130_fd_sc_hd__xnor2_1 _10933_ (.A(_03223_),
    .B(_03231_),
    .Y(_03232_));
 sky130_fd_sc_hd__and2b_1 _10934_ (.A_N(_02504_),
    .B(_02537_),
    .X(_03233_));
 sky130_fd_sc_hd__a21o_1 _10935_ (.A1(_02538_),
    .A2(_02540_),
    .B1(_03233_),
    .X(_03234_));
 sky130_fd_sc_hd__or2_1 _10936_ (.A(_03230_),
    .B(_03229_),
    .X(_03236_));
 sky130_fd_sc_hd__xnor2_2 _10937_ (.A(_03225_),
    .B(_03236_),
    .Y(_03237_));
 sky130_fd_sc_hd__and2b_1 _10938_ (.A_N(_03231_),
    .B(_03223_),
    .X(_03238_));
 sky130_fd_sc_hd__a31o_1 _10939_ (.A1(_03232_),
    .A2(_03234_),
    .A3(_03237_),
    .B1(_03238_),
    .X(_03239_));
 sky130_fd_sc_hd__o21a_1 _10940_ (.A1(_03199_),
    .A2(_03204_),
    .B1(_03192_),
    .X(_03240_));
 sky130_fd_sc_hd__o21a_1 _10941_ (.A1(_03215_),
    .A2(_03219_),
    .B1(_03207_),
    .X(_03241_));
 sky130_fd_sc_hd__a211o_1 _10942_ (.A1(_03221_),
    .A2(_03239_),
    .B1(_03240_),
    .C1(_03241_),
    .X(_03242_));
 sky130_fd_sc_hd__and2_1 _10943_ (.A(_03073_),
    .B(_03100_),
    .X(_03243_));
 sky130_fd_sc_hd__nor2_1 _10944_ (.A(_03101_),
    .B(_03243_),
    .Y(_03244_));
 sky130_fd_sc_hd__or2_1 _10945_ (.A(_03244_),
    .B(_03172_),
    .X(_03245_));
 sky130_fd_sc_hd__o21a_1 _10946_ (.A1(_03172_),
    .A2(_03187_),
    .B1(_03244_),
    .X(_03247_));
 sky130_fd_sc_hd__a41o_1 _10947_ (.A1(_03189_),
    .A2(_03205_),
    .A3(_03242_),
    .A4(_03245_),
    .B1(_03247_),
    .X(_03248_));
 sky130_fd_sc_hd__a311o_1 _10948_ (.A1(_03064_),
    .A2(_03067_),
    .A3(_03104_),
    .B1(_03106_),
    .C1(_03065_),
    .X(_03249_));
 sky130_fd_sc_hd__a21oi_2 _10949_ (.A1(_03108_),
    .A2(_03248_),
    .B1(_03249_),
    .Y(_03250_));
 sky130_fd_sc_hd__and4_1 _10950_ (.A(_00143_),
    .B(_04906_),
    .C(_01508_),
    .D(_01504_),
    .X(_03251_));
 sky130_fd_sc_hd__a22o_1 _10951_ (.A1(_00143_),
    .A2(_01508_),
    .B1(_01505_),
    .B2(_04906_),
    .X(_03252_));
 sky130_fd_sc_hd__or2b_1 _10952_ (.A(_03251_),
    .B_N(_03252_),
    .X(_03253_));
 sky130_fd_sc_hd__nand2_1 _10953_ (.A(_00298_),
    .B(_00608_),
    .Y(_03254_));
 sky130_fd_sc_hd__xnor2_1 _10954_ (.A(_03253_),
    .B(_03254_),
    .Y(_03255_));
 sky130_fd_sc_hd__a22o_1 _10955_ (.A1(_04895_),
    .A2(_01507_),
    .B1(_01504_),
    .B2(_04928_),
    .X(_03256_));
 sky130_fd_sc_hd__and4_1 _10956_ (.A(_04895_),
    .B(_04873_),
    .C(_01507_),
    .D(_01504_),
    .X(_03258_));
 sky130_fd_sc_hd__a31o_1 _10957_ (.A1(_00145_),
    .A2(_00608_),
    .A3(_03256_),
    .B1(_03258_),
    .X(_03259_));
 sky130_fd_sc_hd__or2b_1 _10958_ (.A(_03255_),
    .B_N(_03259_),
    .X(_03260_));
 sky130_fd_sc_hd__a31o_1 _10959_ (.A1(_00859_),
    .A2(_01400_),
    .A3(_03252_),
    .B1(_03251_),
    .X(_03261_));
 sky130_fd_sc_hd__and4_1 _10960_ (.A(_00145_),
    .B(_00310_),
    .C(_02187_),
    .D(_02189_),
    .X(_03262_));
 sky130_fd_sc_hd__a22oi_1 _10961_ (.A1(_00859_),
    .A2(_02188_),
    .B1(_02190_),
    .B2(_01472_),
    .Y(_03263_));
 sky130_fd_sc_hd__nor2_1 _10962_ (.A(_03262_),
    .B(_03263_),
    .Y(_03264_));
 sky130_fd_sc_hd__nand2_1 _10963_ (.A(_03261_),
    .B(_03264_),
    .Y(_03265_));
 sky130_fd_sc_hd__or2_1 _10964_ (.A(_03261_),
    .B(_03264_),
    .X(_03266_));
 sky130_fd_sc_hd__and2_1 _10965_ (.A(_03265_),
    .B(_03266_),
    .X(_03267_));
 sky130_fd_sc_hd__and2b_1 _10966_ (.A_N(_03260_),
    .B(_03267_),
    .X(_03269_));
 sky130_fd_sc_hd__xor2_1 _10967_ (.A(_03260_),
    .B(_03267_),
    .X(_03270_));
 sky130_fd_sc_hd__and4_1 _10968_ (.A(_04862_),
    .B(net4),
    .C(net46),
    .D(_01368_),
    .X(_03271_));
 sky130_fd_sc_hd__inv_2 _10969_ (.A(_03271_),
    .Y(_03272_));
 sky130_fd_sc_hd__a22o_1 _10970_ (.A1(_04862_),
    .A2(_00604_),
    .B1(_01506_),
    .B2(_04873_),
    .X(_03273_));
 sky130_fd_sc_hd__and4_1 _10971_ (.A(_00142_),
    .B(_00457_),
    .C(_03272_),
    .D(_03273_),
    .X(_03274_));
 sky130_fd_sc_hd__a22oi_1 _10972_ (.A1(_00145_),
    .A2(_00460_),
    .B1(_03272_),
    .B2(_03273_),
    .Y(_03275_));
 sky130_fd_sc_hd__nor2_1 _10973_ (.A(_03274_),
    .B(_03275_),
    .Y(_03276_));
 sky130_fd_sc_hd__and4_1 _10974_ (.A(_04917_),
    .B(_04939_),
    .C(_00460_),
    .D(_01400_),
    .X(_03277_));
 sky130_fd_sc_hd__nand2_1 _10975_ (.A(_03276_),
    .B(_03277_),
    .Y(_03278_));
 sky130_fd_sc_hd__and2b_1 _10976_ (.A_N(_03258_),
    .B(_03256_),
    .X(_03280_));
 sky130_fd_sc_hd__nand2_1 _10977_ (.A(_00143_),
    .B(_00607_),
    .Y(_03281_));
 sky130_fd_sc_hd__xnor2_1 _10978_ (.A(_03280_),
    .B(_03281_),
    .Y(_03282_));
 sky130_fd_sc_hd__or2_1 _10979_ (.A(_03271_),
    .B(_03274_),
    .X(_03283_));
 sky130_fd_sc_hd__nand2_1 _10980_ (.A(_00158_),
    .B(_00457_),
    .Y(_03284_));
 sky130_fd_sc_hd__xnor2_1 _10981_ (.A(_03283_),
    .B(_03284_),
    .Y(_03285_));
 sky130_fd_sc_hd__nand2_1 _10982_ (.A(_03282_),
    .B(_03285_),
    .Y(_03286_));
 sky130_fd_sc_hd__or2_1 _10983_ (.A(_03282_),
    .B(_03285_),
    .X(_03287_));
 sky130_fd_sc_hd__nand2_1 _10984_ (.A(_03286_),
    .B(_03287_),
    .Y(_03288_));
 sky130_fd_sc_hd__nor2_1 _10985_ (.A(_03278_),
    .B(_03288_),
    .Y(_03289_));
 sky130_fd_sc_hd__inv_2 _10986_ (.A(_03286_),
    .Y(_03291_));
 sky130_fd_sc_hd__a31o_1 _10987_ (.A1(_00310_),
    .A2(_00459_),
    .A3(_03283_),
    .B1(_03291_),
    .X(_03292_));
 sky130_fd_sc_hd__or2b_1 _10988_ (.A(_03259_),
    .B_N(_03255_),
    .X(_03293_));
 sky130_fd_sc_hd__nand2_1 _10989_ (.A(_03260_),
    .B(_03293_),
    .Y(_03294_));
 sky130_fd_sc_hd__or2b_1 _10990_ (.A(_03292_),
    .B_N(_03294_),
    .X(_03295_));
 sky130_fd_sc_hd__and2b_1 _10991_ (.A_N(_03294_),
    .B(_03292_),
    .X(_03296_));
 sky130_fd_sc_hd__a21oi_1 _10992_ (.A1(_03289_),
    .A2(_03295_),
    .B1(_03296_),
    .Y(_03297_));
 sky130_fd_sc_hd__nor2_1 _10993_ (.A(_03270_),
    .B(_03297_),
    .Y(_03298_));
 sky130_fd_sc_hd__nand2_1 _10994_ (.A(_01473_),
    .B(_02188_),
    .Y(_03299_));
 sky130_fd_sc_hd__and3_1 _10995_ (.A(_02247_),
    .B(_02190_),
    .C(_03299_),
    .X(_03300_));
 sky130_fd_sc_hd__xnor2_1 _10996_ (.A(_03265_),
    .B(_03300_),
    .Y(_03302_));
 sky130_fd_sc_hd__o21a_1 _10997_ (.A1(_03269_),
    .A2(_03298_),
    .B1(_03302_),
    .X(_03303_));
 sky130_fd_sc_hd__nor3_1 _10998_ (.A(_03302_),
    .B(_03269_),
    .C(_03298_),
    .Y(_03304_));
 sky130_fd_sc_hd__nor2_2 _10999_ (.A(_03303_),
    .B(_03304_),
    .Y(_03305_));
 sky130_fd_sc_hd__a22o_1 _11000_ (.A1(_04378_),
    .A2(net47),
    .B1(_00959_),
    .B2(_02971_),
    .X(_03306_));
 sky130_fd_sc_hd__and4_1 _11001_ (.A(_02971_),
    .B(_04378_),
    .C(net47),
    .D(_00959_),
    .X(_03307_));
 sky130_fd_sc_hd__a31oi_2 _11002_ (.A1(_05181_),
    .A2(_00604_),
    .A3(_03306_),
    .B1(_03307_),
    .Y(_03308_));
 sky130_fd_sc_hd__and4_1 _11003_ (.A(_05192_),
    .B(_04598_),
    .C(_01368_),
    .D(_00959_),
    .X(_03309_));
 sky130_fd_sc_hd__a22oi_1 _11004_ (.A1(_04598_),
    .A2(_01506_),
    .B1(_01369_),
    .B2(_05203_),
    .Y(_03310_));
 sky130_fd_sc_hd__or2_1 _11005_ (.A(_03309_),
    .B(_03310_),
    .X(_03311_));
 sky130_fd_sc_hd__nor2_1 _11006_ (.A(_03308_),
    .B(_03311_),
    .Y(_03313_));
 sky130_fd_sc_hd__nand2_1 _11007_ (.A(_00293_),
    .B(_01664_),
    .Y(_03314_));
 sky130_fd_sc_hd__and3_1 _11008_ (.A(_00294_),
    .B(_01505_),
    .C(_03314_),
    .X(_03315_));
 sky130_fd_sc_hd__a32o_1 _11009_ (.A1(_05203_),
    .A2(_00604_),
    .A3(_02549_),
    .B1(_02548_),
    .B2(_01369_),
    .X(_03316_));
 sky130_fd_sc_hd__and2b_1 _11010_ (.A_N(_03307_),
    .B(_03306_),
    .X(_03317_));
 sky130_fd_sc_hd__nand2_1 _11011_ (.A(_04598_),
    .B(_00604_),
    .Y(_03318_));
 sky130_fd_sc_hd__xnor2_1 _11012_ (.A(_03317_),
    .B(_03318_),
    .Y(_03319_));
 sky130_fd_sc_hd__xor2_1 _11013_ (.A(_03308_),
    .B(_03311_),
    .X(_03320_));
 sky130_fd_sc_hd__and3_1 _11014_ (.A(_03316_),
    .B(_03319_),
    .C(_03320_),
    .X(_03321_));
 sky130_fd_sc_hd__and3_1 _11015_ (.A(_05181_),
    .B(net45),
    .C(_02553_),
    .X(_03322_));
 sky130_fd_sc_hd__a21o_1 _11016_ (.A1(_02552_),
    .A2(_02556_),
    .B1(_03322_),
    .X(_03324_));
 sky130_fd_sc_hd__xor2_1 _11017_ (.A(_03316_),
    .B(_03319_),
    .X(_03325_));
 sky130_fd_sc_hd__and2_1 _11018_ (.A(_03324_),
    .B(_03325_),
    .X(_03326_));
 sky130_fd_sc_hd__xnor2_1 _11019_ (.A(_03324_),
    .B(_03325_),
    .Y(_03327_));
 sky130_fd_sc_hd__nor2_1 _11020_ (.A(_02558_),
    .B(_03327_),
    .Y(_03328_));
 sky130_fd_sc_hd__a21oi_1 _11021_ (.A1(_03316_),
    .A2(_03319_),
    .B1(_03320_),
    .Y(_03329_));
 sky130_fd_sc_hd__nor2_1 _11022_ (.A(_03321_),
    .B(_03329_),
    .Y(_03330_));
 sky130_fd_sc_hd__o21a_1 _11023_ (.A1(_03326_),
    .A2(_03328_),
    .B1(_03330_),
    .X(_03331_));
 sky130_fd_sc_hd__xor2_1 _11024_ (.A(_03313_),
    .B(_03315_),
    .X(_03332_));
 sky130_fd_sc_hd__o21a_1 _11025_ (.A1(_03321_),
    .A2(_03331_),
    .B1(_03332_),
    .X(_03333_));
 sky130_fd_sc_hd__a211o_1 _11026_ (.A1(_03313_),
    .A2(_03315_),
    .B1(_03333_),
    .C1(_03309_),
    .X(_03335_));
 sky130_fd_sc_hd__a22o_1 _11027_ (.A1(_05027_),
    .A2(_00780_),
    .B1(_00777_),
    .B2(_04851_),
    .X(_03336_));
 sky130_fd_sc_hd__and4_1 _11028_ (.A(net6),
    .B(_04851_),
    .C(_00780_),
    .D(_00777_),
    .X(_03337_));
 sky130_fd_sc_hd__a31oi_2 _11029_ (.A1(_00158_),
    .A2(_04037_),
    .A3(_03336_),
    .B1(_03337_),
    .Y(_03338_));
 sky130_fd_sc_hd__and4_1 _11030_ (.A(_05027_),
    .B(net7),
    .C(_00612_),
    .D(_00613_),
    .X(_03339_));
 sky130_fd_sc_hd__a22oi_1 _11031_ (.A1(net7),
    .A2(_00782_),
    .B1(_00778_),
    .B2(_05027_),
    .Y(_03340_));
 sky130_fd_sc_hd__or2_1 _11032_ (.A(_03339_),
    .B(_03340_),
    .X(_03341_));
 sky130_fd_sc_hd__nor2_1 _11033_ (.A(_03338_),
    .B(_03341_),
    .Y(_03342_));
 sky130_fd_sc_hd__nand2_1 _11034_ (.A(_00143_),
    .B(_01518_),
    .Y(_03343_));
 sky130_fd_sc_hd__and3_1 _11035_ (.A(_00298_),
    .B(_01517_),
    .C(_03343_),
    .X(_03344_));
 sky130_fd_sc_hd__a32o_1 _11036_ (.A1(_00142_),
    .A2(_04037_),
    .A3(_02566_),
    .B1(_02564_),
    .B2(_00778_),
    .X(_03346_));
 sky130_fd_sc_hd__and2b_1 _11037_ (.A_N(_03337_),
    .B(_03336_),
    .X(_03347_));
 sky130_fd_sc_hd__nand2_1 _11038_ (.A(net7),
    .B(_00373_),
    .Y(_03348_));
 sky130_fd_sc_hd__xnor2_2 _11039_ (.A(_03347_),
    .B(_03348_),
    .Y(_03349_));
 sky130_fd_sc_hd__xor2_1 _11040_ (.A(_03338_),
    .B(_03341_),
    .X(_03350_));
 sky130_fd_sc_hd__and3_1 _11041_ (.A(_03346_),
    .B(_03349_),
    .C(_03350_),
    .X(_03351_));
 sky130_fd_sc_hd__and3_1 _11042_ (.A(_00158_),
    .B(_04059_),
    .C(_02570_),
    .X(_03352_));
 sky130_fd_sc_hd__a21o_1 _11043_ (.A1(_02569_),
    .A2(_02572_),
    .B1(_03352_),
    .X(_03353_));
 sky130_fd_sc_hd__xor2_1 _11044_ (.A(_03346_),
    .B(_03349_),
    .X(_03354_));
 sky130_fd_sc_hd__and2_1 _11045_ (.A(_03353_),
    .B(_03354_),
    .X(_03355_));
 sky130_fd_sc_hd__xnor2_1 _11046_ (.A(_03353_),
    .B(_03354_),
    .Y(_03357_));
 sky130_fd_sc_hd__nor2_1 _11047_ (.A(_02574_),
    .B(_03357_),
    .Y(_03358_));
 sky130_fd_sc_hd__a21oi_1 _11048_ (.A1(_03346_),
    .A2(_03349_),
    .B1(_03350_),
    .Y(_03359_));
 sky130_fd_sc_hd__nor2_1 _11049_ (.A(_03351_),
    .B(_03359_),
    .Y(_03360_));
 sky130_fd_sc_hd__o21a_1 _11050_ (.A1(_03355_),
    .A2(_03358_),
    .B1(_03360_),
    .X(_03361_));
 sky130_fd_sc_hd__xor2_1 _11051_ (.A(_03342_),
    .B(_03344_),
    .X(_03362_));
 sky130_fd_sc_hd__o21a_1 _11052_ (.A1(_03351_),
    .A2(_03361_),
    .B1(_03362_),
    .X(_03363_));
 sky130_fd_sc_hd__a211o_1 _11053_ (.A1(_03342_),
    .A2(_03344_),
    .B1(_03363_),
    .C1(_03339_),
    .X(_03364_));
 sky130_fd_sc_hd__and2_1 _11054_ (.A(_03335_),
    .B(_03364_),
    .X(_03365_));
 sky130_fd_sc_hd__or2b_1 _11055_ (.A(_03296_),
    .B_N(_03295_),
    .X(_03366_));
 sky130_fd_sc_hd__xnor2_1 _11056_ (.A(_03289_),
    .B(_03366_),
    .Y(_03368_));
 sky130_fd_sc_hd__and2_1 _11057_ (.A(_03365_),
    .B(_03368_),
    .X(_03369_));
 sky130_fd_sc_hd__nor2_1 _11058_ (.A(_03365_),
    .B(_03368_),
    .Y(_03370_));
 sky130_fd_sc_hd__or2_1 _11059_ (.A(_03369_),
    .B(_03370_),
    .X(_03371_));
 sky130_fd_sc_hd__and2_1 _11060_ (.A(_03278_),
    .B(_03288_),
    .X(_03372_));
 sky130_fd_sc_hd__nor2_1 _11061_ (.A(_03289_),
    .B(_03372_),
    .Y(_03373_));
 sky130_fd_sc_hd__nor3_1 _11062_ (.A(_03332_),
    .B(_03321_),
    .C(_03331_),
    .Y(_03374_));
 sky130_fd_sc_hd__nor2_1 _11063_ (.A(_03333_),
    .B(_03374_),
    .Y(_03375_));
 sky130_fd_sc_hd__nor3_1 _11064_ (.A(_03362_),
    .B(_03351_),
    .C(_03361_),
    .Y(_03376_));
 sky130_fd_sc_hd__nor2_1 _11065_ (.A(_03363_),
    .B(_03376_),
    .Y(_03377_));
 sky130_fd_sc_hd__nand2_1 _11066_ (.A(_03375_),
    .B(_03377_),
    .Y(_03379_));
 sky130_fd_sc_hd__xnor2_1 _11067_ (.A(_03335_),
    .B(_03364_),
    .Y(_03380_));
 sky130_fd_sc_hd__nand2_1 _11068_ (.A(_03379_),
    .B(_03380_),
    .Y(_03381_));
 sky130_fd_sc_hd__nor2_1 _11069_ (.A(_03379_),
    .B(_03380_),
    .Y(_03382_));
 sky130_fd_sc_hd__a21oi_1 _11070_ (.A1(_03373_),
    .A2(_03381_),
    .B1(_03382_),
    .Y(_03383_));
 sky130_fd_sc_hd__nor2_1 _11071_ (.A(_03371_),
    .B(_03383_),
    .Y(_03384_));
 sky130_fd_sc_hd__and2_1 _11072_ (.A(_03371_),
    .B(_03383_),
    .X(_03385_));
 sky130_fd_sc_hd__nor2_1 _11073_ (.A(_03384_),
    .B(_03385_),
    .Y(_03386_));
 sky130_fd_sc_hd__and2b_1 _11074_ (.A_N(_03382_),
    .B(_03381_),
    .X(_03387_));
 sky130_fd_sc_hd__xor2_1 _11075_ (.A(_03373_),
    .B(_03387_),
    .X(_03388_));
 sky130_fd_sc_hd__nor3_1 _11076_ (.A(_03330_),
    .B(_03326_),
    .C(_03328_),
    .Y(_03390_));
 sky130_fd_sc_hd__nor2_1 _11077_ (.A(_03331_),
    .B(_03390_),
    .Y(_03391_));
 sky130_fd_sc_hd__nor3_1 _11078_ (.A(_03360_),
    .B(_03355_),
    .C(_03358_),
    .Y(_03392_));
 sky130_fd_sc_hd__nor2_1 _11079_ (.A(_03361_),
    .B(_03392_),
    .Y(_03393_));
 sky130_fd_sc_hd__nand2_1 _11080_ (.A(_03391_),
    .B(_03393_),
    .Y(_03394_));
 sky130_fd_sc_hd__xnor2_1 _11081_ (.A(_03375_),
    .B(_03377_),
    .Y(_03395_));
 sky130_fd_sc_hd__nor2_1 _11082_ (.A(_03394_),
    .B(_03395_),
    .Y(_03396_));
 sky130_fd_sc_hd__or2_1 _11083_ (.A(_03276_),
    .B(_03277_),
    .X(_03397_));
 sky130_fd_sc_hd__nand2_2 _11084_ (.A(_03278_),
    .B(_03397_),
    .Y(_03398_));
 sky130_fd_sc_hd__and2_1 _11085_ (.A(_03394_),
    .B(_03395_),
    .X(_03399_));
 sky130_fd_sc_hd__nor2_1 _11086_ (.A(_03398_),
    .B(_03399_),
    .Y(_03401_));
 sky130_fd_sc_hd__or3_2 _11087_ (.A(_03388_),
    .B(_03396_),
    .C(_03401_),
    .X(_03402_));
 sky130_fd_sc_hd__nor2_2 _11088_ (.A(_03396_),
    .B(_03399_),
    .Y(_03403_));
 sky130_fd_sc_hd__xnor2_4 _11089_ (.A(_03398_),
    .B(_03403_),
    .Y(_03404_));
 sky130_fd_sc_hd__and2_1 _11090_ (.A(_02558_),
    .B(_03327_),
    .X(_03405_));
 sky130_fd_sc_hd__nor2_1 _11091_ (.A(_03328_),
    .B(_03405_),
    .Y(_03406_));
 sky130_fd_sc_hd__and2_1 _11092_ (.A(_02574_),
    .B(_03357_),
    .X(_03407_));
 sky130_fd_sc_hd__nor2_1 _11093_ (.A(_03358_),
    .B(_03407_),
    .Y(_03408_));
 sky130_fd_sc_hd__nand2_1 _11094_ (.A(_03406_),
    .B(_03408_),
    .Y(_03409_));
 sky130_fd_sc_hd__xnor2_1 _11095_ (.A(_03391_),
    .B(_03393_),
    .Y(_03410_));
 sky130_fd_sc_hd__nor2_1 _11096_ (.A(_03409_),
    .B(_03410_),
    .Y(_03412_));
 sky130_fd_sc_hd__and2_1 _11097_ (.A(_03409_),
    .B(_03410_),
    .X(_03413_));
 sky130_fd_sc_hd__clkbuf_4 _11098_ (.A(_01400_),
    .X(_03414_));
 sky130_fd_sc_hd__a22oi_1 _11099_ (.A1(_00635_),
    .A2(_01066_),
    .B1(_03414_),
    .B2(_07040_),
    .Y(_03415_));
 sky130_fd_sc_hd__nor2_1 _11100_ (.A(_03277_),
    .B(_03415_),
    .Y(_03416_));
 sky130_fd_sc_hd__and2b_1 _11101_ (.A_N(_03413_),
    .B(_03416_),
    .X(_03417_));
 sky130_fd_sc_hd__nor2_2 _11102_ (.A(_03412_),
    .B(_03417_),
    .Y(_03418_));
 sky130_fd_sc_hd__xnor2_4 _11103_ (.A(_03404_),
    .B(_03418_),
    .Y(_03419_));
 sky130_fd_sc_hd__or2_1 _11104_ (.A(_03412_),
    .B(_03413_),
    .X(_03420_));
 sky130_fd_sc_hd__xnor2_1 _11105_ (.A(_03416_),
    .B(_03420_),
    .Y(_03421_));
 sky130_fd_sc_hd__and2_1 _11106_ (.A(_07040_),
    .B(_01066_),
    .X(_03423_));
 sky130_fd_sc_hd__and2_1 _11107_ (.A(_02562_),
    .B(_02577_),
    .X(_03424_));
 sky130_fd_sc_hd__or2_1 _11108_ (.A(_03406_),
    .B(_03408_),
    .X(_03425_));
 sky130_fd_sc_hd__nand2_1 _11109_ (.A(_03409_),
    .B(_03425_),
    .Y(_03426_));
 sky130_fd_sc_hd__nor3_1 _11110_ (.A(_02561_),
    .B(_03424_),
    .C(_03426_),
    .Y(_03427_));
 sky130_fd_sc_hd__o21a_1 _11111_ (.A1(_02561_),
    .A2(_03424_),
    .B1(_03426_),
    .X(_03428_));
 sky130_fd_sc_hd__o21bai_1 _11112_ (.A1(_03423_),
    .A2(_03427_),
    .B1_N(_03428_),
    .Y(_03429_));
 sky130_fd_sc_hd__xnor2_1 _11113_ (.A(_03421_),
    .B(_03429_),
    .Y(_03430_));
 sky130_fd_sc_hd__or2b_1 _11114_ (.A(_02578_),
    .B_N(_02545_),
    .X(_03431_));
 sky130_fd_sc_hd__and2b_1 _11115_ (.A_N(_02545_),
    .B(_02578_),
    .X(_03432_));
 sky130_fd_sc_hd__a21o_1 _11116_ (.A1(_03431_),
    .A2(_02581_),
    .B1(_03432_),
    .X(_03434_));
 sky130_fd_sc_hd__or2_1 _11117_ (.A(_03428_),
    .B(_03427_),
    .X(_03435_));
 sky130_fd_sc_hd__xnor2_2 _11118_ (.A(_03423_),
    .B(_03435_),
    .Y(_03436_));
 sky130_fd_sc_hd__and2b_1 _11119_ (.A_N(_03429_),
    .B(_03421_),
    .X(_03437_));
 sky130_fd_sc_hd__a31o_2 _11120_ (.A1(_03430_),
    .A2(_03434_),
    .A3(_03436_),
    .B1(_03437_),
    .X(_03438_));
 sky130_fd_sc_hd__o21a_1 _11121_ (.A1(_03396_),
    .A2(_03401_),
    .B1(_03388_),
    .X(_03439_));
 sky130_fd_sc_hd__o21a_1 _11122_ (.A1(_03412_),
    .A2(_03417_),
    .B1(_03404_),
    .X(_03440_));
 sky130_fd_sc_hd__a211o_1 _11123_ (.A1(_03419_),
    .A2(_03438_),
    .B1(_03439_),
    .C1(_03440_),
    .X(_03441_));
 sky130_fd_sc_hd__and2_1 _11124_ (.A(_03270_),
    .B(_03297_),
    .X(_03442_));
 sky130_fd_sc_hd__nor2_1 _11125_ (.A(_03298_),
    .B(_03442_),
    .Y(_03443_));
 sky130_fd_sc_hd__or2_1 _11126_ (.A(_03443_),
    .B(_03369_),
    .X(_03445_));
 sky130_fd_sc_hd__o21a_1 _11127_ (.A1(_03369_),
    .A2(_03384_),
    .B1(_03443_),
    .X(_03446_));
 sky130_fd_sc_hd__a41o_1 _11128_ (.A1(_03386_),
    .A2(_03402_),
    .A3(_03441_),
    .A4(_03445_),
    .B1(_03446_),
    .X(_03447_));
 sky130_fd_sc_hd__a311o_1 _11129_ (.A1(_03261_),
    .A2(_03264_),
    .A3(_03300_),
    .B1(_03303_),
    .C1(_03262_),
    .X(_03448_));
 sky130_fd_sc_hd__a21oi_2 _11130_ (.A1(_03305_),
    .A2(_03447_),
    .B1(_03448_),
    .Y(_03449_));
 sky130_fd_sc_hd__nor2_1 _11131_ (.A(_03250_),
    .B(_03449_),
    .Y(_03450_));
 sky130_fd_sc_hd__or3_1 _11132_ (.A(_03049_),
    .B(_03016_),
    .C(_03045_),
    .X(_03451_));
 sky130_fd_sc_hd__and2_1 _11133_ (.A(_03050_),
    .B(_03451_),
    .X(_03452_));
 sky130_fd_sc_hd__and2_2 _11134_ (.A(_03450_),
    .B(_03452_),
    .X(_03453_));
 sky130_fd_sc_hd__nand2_1 _11135_ (.A(_03002_),
    .B(_03453_),
    .Y(_03454_));
 sky130_fd_sc_hd__nor2_1 _11136_ (.A(_03053_),
    .B(_03454_),
    .Y(_03456_));
 sky130_fd_sc_hd__nor2_1 _11137_ (.A(_03450_),
    .B(_03452_),
    .Y(_03457_));
 sky130_fd_sc_hd__or2_2 _11138_ (.A(_03453_),
    .B(_03457_),
    .X(_03458_));
 sky130_fd_sc_hd__xor2_2 _11139_ (.A(_03108_),
    .B(_03248_),
    .X(_03459_));
 sky130_fd_sc_hd__xor2_2 _11140_ (.A(_03305_),
    .B(_03447_),
    .X(_03460_));
 sky130_fd_sc_hd__and2_2 _11141_ (.A(_03459_),
    .B(_03460_),
    .X(_03461_));
 sky130_fd_sc_hd__xor2_2 _11142_ (.A(_03250_),
    .B(_03449_),
    .X(_03462_));
 sky130_fd_sc_hd__nor3_1 _11143_ (.A(_03044_),
    .B(_03029_),
    .C(_03042_),
    .Y(_03463_));
 sky130_fd_sc_hd__nor2_2 _11144_ (.A(_03045_),
    .B(_03463_),
    .Y(_03464_));
 sky130_fd_sc_hd__a21o_1 _11145_ (.A1(_03461_),
    .A2(_03462_),
    .B1(_03464_),
    .X(_03465_));
 sky130_fd_sc_hd__o21ai_2 _11146_ (.A1(_03461_),
    .A2(_03462_),
    .B1(_03465_),
    .Y(_03467_));
 sky130_fd_sc_hd__nor2_1 _11147_ (.A(_03458_),
    .B(_03467_),
    .Y(_03468_));
 sky130_fd_sc_hd__o21a_1 _11148_ (.A1(_03038_),
    .A2(_03040_),
    .B1(_03031_),
    .X(_03469_));
 sky130_fd_sc_hd__nor2_2 _11149_ (.A(_03042_),
    .B(_03469_),
    .Y(_03470_));
 sky130_fd_sc_hd__xnor2_2 _11150_ (.A(_03459_),
    .B(_03460_),
    .Y(_03471_));
 sky130_fd_sc_hd__nand2_1 _11151_ (.A(_03244_),
    .B(_03172_),
    .Y(_03472_));
 sky130_fd_sc_hd__nand2_1 _11152_ (.A(_03245_),
    .B(_03472_),
    .Y(_03473_));
 sky130_fd_sc_hd__a31o_1 _11153_ (.A1(_03189_),
    .A2(_03205_),
    .A3(_03242_),
    .B1(_03187_),
    .X(_03474_));
 sky130_fd_sc_hd__xnor2_2 _11154_ (.A(_03473_),
    .B(_03474_),
    .Y(_03475_));
 sky130_fd_sc_hd__nand2_1 _11155_ (.A(_03443_),
    .B(_03369_),
    .Y(_03476_));
 sky130_fd_sc_hd__nand2_2 _11156_ (.A(_03445_),
    .B(_03476_),
    .Y(_03478_));
 sky130_fd_sc_hd__a31o_2 _11157_ (.A1(_03386_),
    .A2(_03402_),
    .A3(_03441_),
    .B1(_03384_),
    .X(_03479_));
 sky130_fd_sc_hd__xnor2_4 _11158_ (.A(_03478_),
    .B(_03479_),
    .Y(_03480_));
 sky130_fd_sc_hd__nand2_2 _11159_ (.A(_03475_),
    .B(_03480_),
    .Y(_03481_));
 sky130_fd_sc_hd__nand2_1 _11160_ (.A(_03471_),
    .B(_03481_),
    .Y(_03482_));
 sky130_fd_sc_hd__nor2_1 _11161_ (.A(_03471_),
    .B(_03481_),
    .Y(_03483_));
 sky130_fd_sc_hd__a21o_2 _11162_ (.A1(_03470_),
    .A2(_03482_),
    .B1(_03483_),
    .X(_03484_));
 sky130_fd_sc_hd__xnor2_2 _11163_ (.A(_03461_),
    .B(_03462_),
    .Y(_03485_));
 sky130_fd_sc_hd__xnor2_4 _11164_ (.A(_03464_),
    .B(_03485_),
    .Y(_03486_));
 sky130_fd_sc_hd__and2_1 _11165_ (.A(_03484_),
    .B(_03486_),
    .X(_03487_));
 sky130_fd_sc_hd__nand2_1 _11166_ (.A(_03458_),
    .B(_03467_),
    .Y(_03489_));
 sky130_fd_sc_hd__o21a_1 _11167_ (.A1(_03468_),
    .A2(_03487_),
    .B1(_03489_),
    .X(_03490_));
 sky130_fd_sc_hd__and2_1 _11168_ (.A(_03003_),
    .B(_03050_),
    .X(_03491_));
 sky130_fd_sc_hd__nor2_1 _11169_ (.A(_03051_),
    .B(_03491_),
    .Y(_03492_));
 sky130_fd_sc_hd__o21ai_4 _11170_ (.A1(_03453_),
    .A2(_03492_),
    .B1(_03454_),
    .Y(_03493_));
 sky130_fd_sc_hd__or2_1 _11171_ (.A(_03053_),
    .B(_03493_),
    .X(_03494_));
 sky130_fd_sc_hd__inv_2 _11172_ (.A(_03494_),
    .Y(_03495_));
 sky130_fd_sc_hd__and2_1 _11173_ (.A(_03490_),
    .B(_03495_),
    .X(_03496_));
 sky130_fd_sc_hd__xnor2_2 _11174_ (.A(_03471_),
    .B(_03481_),
    .Y(_03497_));
 sky130_fd_sc_hd__xnor2_4 _11175_ (.A(_03470_),
    .B(_03497_),
    .Y(_03498_));
 sky130_fd_sc_hd__and3_1 _11176_ (.A(_03189_),
    .B(_03205_),
    .C(_03242_),
    .X(_03500_));
 sky130_fd_sc_hd__and3_1 _11177_ (.A(_03386_),
    .B(_03402_),
    .C(_03441_),
    .X(_03501_));
 sky130_fd_sc_hd__a21oi_1 _11178_ (.A1(_03205_),
    .A2(_03242_),
    .B1(_03189_),
    .Y(_03502_));
 sky130_fd_sc_hd__a21oi_2 _11179_ (.A1(_03402_),
    .A2(_03441_),
    .B1(_03386_),
    .Y(_03503_));
 sky130_fd_sc_hd__nor4_1 _11180_ (.A(_03500_),
    .B(_03501_),
    .C(_03502_),
    .D(_03503_),
    .Y(_03504_));
 sky130_fd_sc_hd__xor2_2 _11181_ (.A(_03475_),
    .B(_03480_),
    .X(_03505_));
 sky130_fd_sc_hd__nor2_1 _11182_ (.A(net138),
    .B(_03505_),
    .Y(_03506_));
 sky130_fd_sc_hd__and2_1 _11183_ (.A(_03038_),
    .B(_03040_),
    .X(_03507_));
 sky130_fd_sc_hd__nor2_1 _11184_ (.A(_03041_),
    .B(_03507_),
    .Y(_03508_));
 sky130_fd_sc_hd__a21o_1 _11185_ (.A1(net138),
    .A2(_03505_),
    .B1(_03508_),
    .X(_03509_));
 sky130_fd_sc_hd__and2b_2 _11186_ (.A_N(_03506_),
    .B(_03509_),
    .X(_03511_));
 sky130_fd_sc_hd__and2_1 _11187_ (.A(_03498_),
    .B(_03511_),
    .X(_03512_));
 sky130_fd_sc_hd__xnor2_1 _11188_ (.A(net138),
    .B(_03505_),
    .Y(_03513_));
 sky130_fd_sc_hd__o2bb2a_1 _11189_ (.A1_N(_03508_),
    .A2_N(_03513_),
    .B1(_03509_),
    .B2(_03506_),
    .X(_03514_));
 sky130_fd_sc_hd__inv_2 _11190_ (.A(_03034_),
    .Y(_03515_));
 sky130_fd_sc_hd__o211ai_1 _11191_ (.A1(_03515_),
    .A2(_03035_),
    .B1(_01156_),
    .C1(_01108_),
    .Y(_03516_));
 sky130_fd_sc_hd__a211o_1 _11192_ (.A1(_01156_),
    .A2(_01108_),
    .B1(_03515_),
    .C1(_03035_),
    .X(_03517_));
 sky130_fd_sc_hd__nand2_1 _11193_ (.A(_03516_),
    .B(_03517_),
    .Y(_03518_));
 sky130_fd_sc_hd__a21oi_1 _11194_ (.A1(_03221_),
    .A2(_03239_),
    .B1(_03241_),
    .Y(_03519_));
 sky130_fd_sc_hd__nor3_1 _11195_ (.A(_03192_),
    .B(_03199_),
    .C(_03204_),
    .Y(_03520_));
 sky130_fd_sc_hd__nor2_1 _11196_ (.A(_03520_),
    .B(_03240_),
    .Y(_03522_));
 sky130_fd_sc_hd__xnor2_2 _11197_ (.A(_03519_),
    .B(_03522_),
    .Y(_03523_));
 sky130_fd_sc_hd__a21oi_2 _11198_ (.A1(_03419_),
    .A2(_03438_),
    .B1(_03440_),
    .Y(_03524_));
 sky130_fd_sc_hd__nor3_1 _11199_ (.A(_03388_),
    .B(_03396_),
    .C(_03401_),
    .Y(_03525_));
 sky130_fd_sc_hd__nor2_2 _11200_ (.A(_03525_),
    .B(_03439_),
    .Y(_03526_));
 sky130_fd_sc_hd__xnor2_4 _11201_ (.A(_03524_),
    .B(_03526_),
    .Y(_03527_));
 sky130_fd_sc_hd__nand2_1 _11202_ (.A(_03523_),
    .B(_03527_),
    .Y(_03528_));
 sky130_fd_sc_hd__o22a_1 _11203_ (.A1(_03500_),
    .A2(_03502_),
    .B1(_03503_),
    .B2(_03501_),
    .X(_03529_));
 sky130_fd_sc_hd__nor3_1 _11204_ (.A(net178),
    .B(_03528_),
    .C(_03529_),
    .Y(_03530_));
 sky130_fd_sc_hd__o21a_1 _11205_ (.A1(net178),
    .A2(_03529_),
    .B1(_03528_),
    .X(_03531_));
 sky130_fd_sc_hd__o21ba_1 _11206_ (.A1(_03518_),
    .A2(_03530_),
    .B1_N(_03531_),
    .X(_03533_));
 sky130_fd_sc_hd__and2b_1 _11207_ (.A_N(_03514_),
    .B(_03533_),
    .X(_03534_));
 sky130_fd_sc_hd__or2_1 _11208_ (.A(_03498_),
    .B(_03511_),
    .X(_03535_));
 sky130_fd_sc_hd__o21a_1 _11209_ (.A1(_03512_),
    .A2(_03534_),
    .B1(_03535_),
    .X(_03536_));
 sky130_fd_sc_hd__nor2_1 _11210_ (.A(_02502_),
    .B(_02541_),
    .Y(_03537_));
 sky130_fd_sc_hd__a21oi_2 _11211_ (.A1(_02502_),
    .A2(_02541_),
    .B1(_02582_),
    .Y(_03538_));
 sky130_fd_sc_hd__xor2_1 _11212_ (.A(_03234_),
    .B(_03237_),
    .X(_03539_));
 sky130_fd_sc_hd__xor2_2 _11213_ (.A(_03434_),
    .B(_03436_),
    .X(_03540_));
 sky130_fd_sc_hd__and2_1 _11214_ (.A(_03539_),
    .B(_03540_),
    .X(_03541_));
 sky130_fd_sc_hd__nor2_1 _11215_ (.A(_03539_),
    .B(_03540_),
    .Y(_03542_));
 sky130_fd_sc_hd__or2_1 _11216_ (.A(_03541_),
    .B(_03542_),
    .X(_03544_));
 sky130_fd_sc_hd__o21ai_2 _11217_ (.A1(_03537_),
    .A2(_03538_),
    .B1(_03544_),
    .Y(_03545_));
 sky130_fd_sc_hd__or3_1 _11218_ (.A(_03537_),
    .B(_03544_),
    .C(_03538_),
    .X(_03546_));
 sky130_fd_sc_hd__nand2_2 _11219_ (.A(_00410_),
    .B(_01108_),
    .Y(_03547_));
 sky130_fd_sc_hd__a21o_1 _11220_ (.A1(_03545_),
    .A2(_03546_),
    .B1(_03547_),
    .X(_03548_));
 sky130_fd_sc_hd__nand3_2 _11221_ (.A(_03545_),
    .B(_03547_),
    .C(_03546_),
    .Y(_03549_));
 sky130_fd_sc_hd__nand2_1 _11222_ (.A(_02583_),
    .B(_02586_),
    .Y(_03550_));
 sky130_fd_sc_hd__a21o_1 _11223_ (.A1(_03548_),
    .A2(_03549_),
    .B1(_03550_),
    .X(_03551_));
 sky130_fd_sc_hd__a211o_1 _11224_ (.A1(_03548_),
    .A2(_03549_),
    .B1(_02382_),
    .C1(_02588_),
    .X(_03552_));
 sky130_fd_sc_hd__and3_1 _11225_ (.A(_03232_),
    .B(_03234_),
    .C(_03237_),
    .X(_03553_));
 sky130_fd_sc_hd__a21oi_1 _11226_ (.A1(_03234_),
    .A2(_03237_),
    .B1(_03232_),
    .Y(_03555_));
 sky130_fd_sc_hd__or2_1 _11227_ (.A(_03553_),
    .B(_03555_),
    .X(_03556_));
 sky130_fd_sc_hd__and3_1 _11228_ (.A(_03430_),
    .B(_03434_),
    .C(_03436_),
    .X(_03557_));
 sky130_fd_sc_hd__a21oi_1 _11229_ (.A1(_03434_),
    .A2(_03436_),
    .B1(_03430_),
    .Y(_03558_));
 sky130_fd_sc_hd__or2_1 _11230_ (.A(_03557_),
    .B(_03558_),
    .X(_03559_));
 sky130_fd_sc_hd__or2_2 _11231_ (.A(_03556_),
    .B(_03559_),
    .X(_03560_));
 sky130_fd_sc_hd__nand2_1 _11232_ (.A(_03556_),
    .B(_03559_),
    .Y(_03561_));
 sky130_fd_sc_hd__and3_1 _11233_ (.A(_03560_),
    .B(_03541_),
    .C(_03561_),
    .X(_03562_));
 sky130_fd_sc_hd__a21oi_1 _11234_ (.A1(_03560_),
    .A2(_03561_),
    .B1(_03541_),
    .Y(_03563_));
 sky130_fd_sc_hd__a22oi_1 _11235_ (.A1(_03015_),
    .A2(_01062_),
    .B1(_01415_),
    .B2(_00410_),
    .Y(_03564_));
 sky130_fd_sc_hd__nor2_1 _11236_ (.A(_02979_),
    .B(_03564_),
    .Y(_03566_));
 sky130_fd_sc_hd__and2b_1 _11237_ (.A_N(_03563_),
    .B(_03566_),
    .X(_03567_));
 sky130_fd_sc_hd__or2_1 _11238_ (.A(_02978_),
    .B(_02979_),
    .X(_03568_));
 sky130_fd_sc_hd__nand2_1 _11239_ (.A(_02980_),
    .B(_03568_),
    .Y(_03569_));
 sky130_fd_sc_hd__xor2_2 _11240_ (.A(_03221_),
    .B(_03239_),
    .X(_03570_));
 sky130_fd_sc_hd__xor2_4 _11241_ (.A(_03419_),
    .B(_03438_),
    .X(_03571_));
 sky130_fd_sc_hd__xnor2_2 _11242_ (.A(_03570_),
    .B(_03571_),
    .Y(_03572_));
 sky130_fd_sc_hd__xor2_1 _11243_ (.A(_03572_),
    .B(_03560_),
    .X(_03573_));
 sky130_fd_sc_hd__xnor2_1 _11244_ (.A(_03569_),
    .B(_03573_),
    .Y(_03574_));
 sky130_fd_sc_hd__o21a_1 _11245_ (.A1(_03562_),
    .A2(_03567_),
    .B1(_03574_),
    .X(_03575_));
 sky130_fd_sc_hd__nor3_1 _11246_ (.A(_03574_),
    .B(_03562_),
    .C(_03567_),
    .Y(_03577_));
 sky130_fd_sc_hd__or2_1 _11247_ (.A(_03575_),
    .B(_03577_),
    .X(_03578_));
 sky130_fd_sc_hd__nor2_1 _11248_ (.A(_03562_),
    .B(_03563_),
    .Y(_03579_));
 sky130_fd_sc_hd__xor2_1 _11249_ (.A(_03566_),
    .B(_03579_),
    .X(_03580_));
 sky130_fd_sc_hd__o31ai_2 _11250_ (.A1(_03537_),
    .A2(_03544_),
    .A3(_03538_),
    .B1(_03547_),
    .Y(_03581_));
 sky130_fd_sc_hd__and3_1 _11251_ (.A(_03580_),
    .B(_03545_),
    .C(_03581_),
    .X(_03582_));
 sky130_fd_sc_hd__a21oi_1 _11252_ (.A1(_03545_),
    .A2(_03581_),
    .B1(_03580_),
    .Y(_03583_));
 sky130_fd_sc_hd__or3_1 _11253_ (.A(_03578_),
    .B(_03582_),
    .C(_03583_),
    .X(_03584_));
 sky130_fd_sc_hd__a21o_1 _11254_ (.A1(_03551_),
    .A2(_03552_),
    .B1(_03584_),
    .X(_03585_));
 sky130_fd_sc_hd__a21o_1 _11255_ (.A1(_03548_),
    .A2(_03549_),
    .B1(_02588_),
    .X(_03586_));
 sky130_fd_sc_hd__a2111o_1 _11256_ (.A1(_02299_),
    .A2(_02241_),
    .B1(_02384_),
    .C1(_03586_),
    .D1(_03584_),
    .X(_03588_));
 sky130_fd_sc_hd__nand3_1 _11257_ (.A(_03580_),
    .B(_03545_),
    .C(_03581_),
    .Y(_03589_));
 sky130_fd_sc_hd__o21ba_1 _11258_ (.A1(_03577_),
    .A2(_03589_),
    .B1_N(_03575_),
    .X(_03590_));
 sky130_fd_sc_hd__nand2_1 _11259_ (.A(_03570_),
    .B(_03571_),
    .Y(_03591_));
 sky130_fd_sc_hd__xnor2_2 _11260_ (.A(_03523_),
    .B(_03527_),
    .Y(_03592_));
 sky130_fd_sc_hd__nor2_1 _11261_ (.A(_03591_),
    .B(_03592_),
    .Y(_03593_));
 sky130_fd_sc_hd__and2_1 _11262_ (.A(_02980_),
    .B(_02983_),
    .X(_03594_));
 sky130_fd_sc_hd__nor2_1 _11263_ (.A(_03032_),
    .B(_03594_),
    .Y(_03595_));
 sky130_fd_sc_hd__nand2_1 _11264_ (.A(_03591_),
    .B(_03592_),
    .Y(_03596_));
 sky130_fd_sc_hd__o21ai_2 _11265_ (.A1(_03593_),
    .A2(_03595_),
    .B1(_03596_),
    .Y(_03597_));
 sky130_fd_sc_hd__or3_1 _11266_ (.A(_03531_),
    .B(_03518_),
    .C(_03530_),
    .X(_03599_));
 sky130_fd_sc_hd__o21ai_1 _11267_ (.A1(_03531_),
    .A2(_03530_),
    .B1(_03518_),
    .Y(_03600_));
 sky130_fd_sc_hd__and2_1 _11268_ (.A(_03599_),
    .B(_03600_),
    .X(_03601_));
 sky130_fd_sc_hd__xor2_2 _11269_ (.A(_03597_),
    .B(_03601_),
    .X(_03602_));
 sky130_fd_sc_hd__xnor2_1 _11270_ (.A(_03591_),
    .B(_03592_),
    .Y(_03603_));
 sky130_fd_sc_hd__xnor2_1 _11271_ (.A(_03595_),
    .B(_03603_),
    .Y(_03604_));
 sky130_fd_sc_hd__a21o_1 _11272_ (.A1(_03572_),
    .A2(_03560_),
    .B1(_03569_),
    .X(_03605_));
 sky130_fd_sc_hd__o21a_1 _11273_ (.A1(_03572_),
    .A2(_03560_),
    .B1(_03605_),
    .X(_03606_));
 sky130_fd_sc_hd__inv_2 _11274_ (.A(_03606_),
    .Y(_03607_));
 sky130_fd_sc_hd__and2_1 _11275_ (.A(_03604_),
    .B(_03607_),
    .X(_03608_));
 sky130_fd_sc_hd__or2_1 _11276_ (.A(_03604_),
    .B(_03607_),
    .X(_03610_));
 sky130_fd_sc_hd__and2b_2 _11277_ (.A_N(_03608_),
    .B(_03610_),
    .X(_03611_));
 sky130_fd_sc_hd__nand2_1 _11278_ (.A(_03602_),
    .B(_03611_),
    .Y(_03612_));
 sky130_fd_sc_hd__xor2_4 _11279_ (.A(_03498_),
    .B(_03511_),
    .X(_03613_));
 sky130_fd_sc_hd__xnor2_2 _11280_ (.A(_03514_),
    .B(_03533_),
    .Y(_03614_));
 sky130_fd_sc_hd__nand2_1 _11281_ (.A(_03613_),
    .B(_03614_),
    .Y(_03615_));
 sky130_fd_sc_hd__a311oi_2 _11282_ (.A1(_03585_),
    .A2(_03588_),
    .A3(_03590_),
    .B1(_03612_),
    .C1(_03615_),
    .Y(_03616_));
 sky130_fd_sc_hd__nor2_1 _11283_ (.A(_03597_),
    .B(_03601_),
    .Y(_03617_));
 sky130_fd_sc_hd__nand2_1 _11284_ (.A(_03597_),
    .B(_03601_),
    .Y(_03618_));
 sky130_fd_sc_hd__o21ai_1 _11285_ (.A1(_03617_),
    .A2(_03608_),
    .B1(_03618_),
    .Y(_03619_));
 sky130_fd_sc_hd__nor2_1 _11286_ (.A(_03619_),
    .B(_03615_),
    .Y(_03621_));
 sky130_fd_sc_hd__xor2_2 _11287_ (.A(_03458_),
    .B(_03467_),
    .X(_03622_));
 sky130_fd_sc_hd__xor2_4 _11288_ (.A(_03484_),
    .B(_03486_),
    .X(_03623_));
 sky130_fd_sc_hd__and2_1 _11289_ (.A(_03622_),
    .B(_03623_),
    .X(_03624_));
 sky130_fd_sc_hd__o311a_1 _11290_ (.A1(_03536_),
    .A2(_03616_),
    .A3(_03621_),
    .B1(_03624_),
    .C1(_03495_),
    .X(_03625_));
 sky130_fd_sc_hd__or3_2 _11291_ (.A(_03456_),
    .B(_03496_),
    .C(_03625_),
    .X(_03626_));
 sky130_fd_sc_hd__xnor2_2 _11292_ (.A(_02746_),
    .B(_02790_),
    .Y(_03627_));
 sky130_fd_sc_hd__and2_1 _11293_ (.A(_02757_),
    .B(_02788_),
    .X(_03628_));
 sky130_fd_sc_hd__nor2_1 _11294_ (.A(_02789_),
    .B(_03628_),
    .Y(_03629_));
 sky130_fd_sc_hd__a21bo_1 _11295_ (.A1(_02862_),
    .A2(_02908_),
    .B1_N(_02859_),
    .X(_03630_));
 sky130_fd_sc_hd__and4_1 _11296_ (.A(_00819_),
    .B(_00818_),
    .C(_02736_),
    .D(_02737_),
    .X(_03632_));
 sky130_fd_sc_hd__a211o_1 _11297_ (.A1(_02810_),
    .A2(_02899_),
    .B1(_02901_),
    .C1(_03632_),
    .X(_03633_));
 sky130_fd_sc_hd__o21a_1 _11298_ (.A1(_02910_),
    .A2(_03630_),
    .B1(_03633_),
    .X(_03634_));
 sky130_fd_sc_hd__nor2_1 _11299_ (.A(_02770_),
    .B(_02787_),
    .Y(_03635_));
 sky130_fd_sc_hd__xnor2_1 _11300_ (.A(_02785_),
    .B(_03635_),
    .Y(_03636_));
 sky130_fd_sc_hd__and2_1 _11301_ (.A(_03634_),
    .B(_03636_),
    .X(_03637_));
 sky130_fd_sc_hd__nand2_1 _11302_ (.A(_03629_),
    .B(_03637_),
    .Y(_03638_));
 sky130_fd_sc_hd__or2_1 _11303_ (.A(_03629_),
    .B(_03637_),
    .X(_03639_));
 sky130_fd_sc_hd__and2_1 _11304_ (.A(_03638_),
    .B(_03639_),
    .X(_03640_));
 sky130_fd_sc_hd__nor2_1 _11305_ (.A(_03634_),
    .B(_03636_),
    .Y(_03641_));
 sky130_fd_sc_hd__or2_1 _11306_ (.A(_03637_),
    .B(_03641_),
    .X(_03643_));
 sky130_fd_sc_hd__nor3_1 _11307_ (.A(_02910_),
    .B(_03633_),
    .C(_03630_),
    .Y(_03644_));
 sky130_fd_sc_hd__or2_1 _11308_ (.A(_03634_),
    .B(_03644_),
    .X(_03645_));
 sky130_fd_sc_hd__nand2_1 _11309_ (.A(_02913_),
    .B(_03645_),
    .Y(_03646_));
 sky130_fd_sc_hd__and2_1 _11310_ (.A(_02770_),
    .B(_02787_),
    .X(_03647_));
 sky130_fd_sc_hd__nor2_1 _11311_ (.A(_03635_),
    .B(_03647_),
    .Y(_03648_));
 sky130_fd_sc_hd__nor2_1 _11312_ (.A(_02913_),
    .B(_03645_),
    .Y(_03649_));
 sky130_fd_sc_hd__a21oi_1 _11313_ (.A1(_03646_),
    .A2(_03648_),
    .B1(_03649_),
    .Y(_03650_));
 sky130_fd_sc_hd__or2_1 _11314_ (.A(_03643_),
    .B(_03650_),
    .X(_03651_));
 sky130_fd_sc_hd__nand2_1 _11315_ (.A(_03643_),
    .B(_03650_),
    .Y(_03652_));
 sky130_fd_sc_hd__nand2_1 _11316_ (.A(_03651_),
    .B(_03652_),
    .Y(_03654_));
 sky130_fd_sc_hd__nor2_1 _11317_ (.A(_02796_),
    .B(_02918_),
    .Y(_03655_));
 sky130_fd_sc_hd__or2b_1 _11318_ (.A(_03649_),
    .B_N(_03646_),
    .X(_03656_));
 sky130_fd_sc_hd__xnor2_1 _11319_ (.A(_03648_),
    .B(_03656_),
    .Y(_03657_));
 sky130_fd_sc_hd__o21ai_1 _11320_ (.A1(_02917_),
    .A2(_03655_),
    .B1(_03657_),
    .Y(_03658_));
 sky130_fd_sc_hd__and2_1 _11321_ (.A(_02920_),
    .B(_02932_),
    .X(_03659_));
 sky130_fd_sc_hd__a21oi_2 _11322_ (.A1(_02933_),
    .A2(_03052_),
    .B1(_03659_),
    .Y(_03660_));
 sky130_fd_sc_hd__or3_1 _11323_ (.A(_02917_),
    .B(_03657_),
    .C(_03655_),
    .X(_03661_));
 sky130_fd_sc_hd__a21bo_1 _11324_ (.A1(_03658_),
    .A2(_03660_),
    .B1_N(_03661_),
    .X(_03662_));
 sky130_fd_sc_hd__o21ai_2 _11325_ (.A1(_03654_),
    .A2(_03662_),
    .B1(_03651_),
    .Y(_03663_));
 sky130_fd_sc_hd__nand2_1 _11326_ (.A(_03640_),
    .B(_03663_),
    .Y(_03665_));
 sky130_fd_sc_hd__nand2_1 _11327_ (.A(_03638_),
    .B(_03665_),
    .Y(_03666_));
 sky130_fd_sc_hd__xnor2_2 _11328_ (.A(_03627_),
    .B(_03666_),
    .Y(_03667_));
 sky130_fd_sc_hd__xnor2_2 _11329_ (.A(_03640_),
    .B(_03663_),
    .Y(_03668_));
 sky130_fd_sc_hd__xor2_2 _11330_ (.A(_03654_),
    .B(_03662_),
    .X(_03669_));
 sky130_fd_sc_hd__and2_1 _11331_ (.A(_03661_),
    .B(_03658_),
    .X(_03670_));
 sky130_fd_sc_hd__xnor2_2 _11332_ (.A(_03660_),
    .B(_03670_),
    .Y(_03671_));
 sky130_fd_sc_hd__nand2_1 _11333_ (.A(_03669_),
    .B(_03671_),
    .Y(_03672_));
 sky130_fd_sc_hd__or2_1 _11334_ (.A(_03668_),
    .B(_03672_),
    .X(_03673_));
 sky130_fd_sc_hd__inv_2 _11335_ (.A(_03673_),
    .Y(_03674_));
 sky130_fd_sc_hd__and3_1 _11336_ (.A(_03626_),
    .B(_03667_),
    .C(_03674_),
    .X(_03675_));
 sky130_fd_sc_hd__a21o_1 _11337_ (.A1(_03638_),
    .A2(_03665_),
    .B1(_03627_),
    .X(_03676_));
 sky130_fd_sc_hd__or3b_1 _11338_ (.A(_02793_),
    .B(_03675_),
    .C_N(_03676_),
    .X(_03677_));
 sky130_fd_sc_hd__clkbuf_4 _11339_ (.A(_02673_),
    .X(_03678_));
 sky130_fd_sc_hd__clkbuf_4 _11340_ (.A(_03678_),
    .X(_03679_));
 sky130_fd_sc_hd__clkbuf_4 _11341_ (.A(_03679_),
    .X(_03680_));
 sky130_fd_sc_hd__clkbuf_4 _11342_ (.A(_02459_),
    .X(_03681_));
 sky130_fd_sc_hd__clkbuf_4 _11343_ (.A(_03681_),
    .X(_03682_));
 sky130_fd_sc_hd__clkbuf_4 _11344_ (.A(_03682_),
    .X(_03683_));
 sky130_fd_sc_hd__buf_2 _11345_ (.A(_03683_),
    .X(_03684_));
 sky130_fd_sc_hd__clkbuf_4 _11346_ (.A(_02135_),
    .X(_03686_));
 sky130_fd_sc_hd__clkbuf_4 _11347_ (.A(_03686_),
    .X(_03687_));
 sky130_fd_sc_hd__a22o_1 _11348_ (.A1(_02249_),
    .A2(_01956_),
    .B1(_03687_),
    .B2(_01312_),
    .X(_03688_));
 sky130_fd_sc_hd__and3_1 _11349_ (.A(_02249_),
    .B(_01312_),
    .C(_01956_),
    .X(_03689_));
 sky130_fd_sc_hd__buf_2 _11350_ (.A(_03687_),
    .X(_03690_));
 sky130_fd_sc_hd__a32o_1 _11351_ (.A1(_00544_),
    .A2(_03684_),
    .A3(_03688_),
    .B1(_03689_),
    .B2(_03690_),
    .X(_03691_));
 sky130_fd_sc_hd__and3_1 _11352_ (.A(_01155_),
    .B(_03680_),
    .C(_03691_),
    .X(_03692_));
 sky130_fd_sc_hd__and4_1 _11353_ (.A(_02246_),
    .B(_02249_),
    .C(_01956_),
    .D(_03687_),
    .X(_03693_));
 sky130_fd_sc_hd__a22oi_1 _11354_ (.A1(_02246_),
    .A2(_01957_),
    .B1(_03690_),
    .B2(_02249_),
    .Y(_03694_));
 sky130_fd_sc_hd__and4bb_1 _11355_ (.A_N(_03693_),
    .B_N(_03694_),
    .C(_01312_),
    .D(_03684_),
    .X(_03695_));
 sky130_fd_sc_hd__clkbuf_4 _11356_ (.A(_03684_),
    .X(_03697_));
 sky130_fd_sc_hd__o2bb2a_1 _11357_ (.A1_N(_01312_),
    .A2_N(_03697_),
    .B1(_03693_),
    .B2(_03694_),
    .X(_03698_));
 sky130_fd_sc_hd__clkbuf_4 _11358_ (.A(_03680_),
    .X(_03699_));
 sky130_fd_sc_hd__a21oi_1 _11359_ (.A1(_01155_),
    .A2(_03699_),
    .B1(_03691_),
    .Y(_03700_));
 sky130_fd_sc_hd__nor4_1 _11360_ (.A(_03695_),
    .B(_03692_),
    .C(_03698_),
    .D(_03700_),
    .Y(_03701_));
 sky130_fd_sc_hd__and4_1 _11361_ (.A(_00843_),
    .B(_00844_),
    .C(_03687_),
    .D(_03684_),
    .X(_03702_));
 sky130_fd_sc_hd__a22o_1 _11362_ (.A1(_02246_),
    .A2(_03687_),
    .B1(_03684_),
    .B2(_02249_),
    .X(_03703_));
 sky130_fd_sc_hd__and2b_1 _11363_ (.A_N(_03702_),
    .B(_03703_),
    .X(_03704_));
 sky130_fd_sc_hd__nand2_1 _11364_ (.A(_01312_),
    .B(_03680_),
    .Y(_03705_));
 sky130_fd_sc_hd__xnor2_1 _11365_ (.A(_03704_),
    .B(_03705_),
    .Y(_03706_));
 sky130_fd_sc_hd__o21a_1 _11366_ (.A1(_03693_),
    .A2(_03695_),
    .B1(_03706_),
    .X(_03708_));
 sky130_fd_sc_hd__nor3_1 _11367_ (.A(_03693_),
    .B(_03695_),
    .C(_03706_),
    .Y(_03709_));
 sky130_fd_sc_hd__nor2_1 _11368_ (.A(_03708_),
    .B(_03709_),
    .Y(_03710_));
 sky130_fd_sc_hd__o21a_1 _11369_ (.A1(_03692_),
    .A2(net142),
    .B1(_03710_),
    .X(_03711_));
 sky130_fd_sc_hd__nor3_1 _11370_ (.A(_03692_),
    .B(net142),
    .C(_03710_),
    .Y(_03712_));
 sky130_fd_sc_hd__a21bo_1 _11371_ (.A1(_03690_),
    .A2(_03689_),
    .B1_N(_03688_),
    .X(_03713_));
 sky130_fd_sc_hd__nand2_2 _11372_ (.A(_01155_),
    .B(_03697_),
    .Y(_03714_));
 sky130_fd_sc_hd__xnor2_4 _11373_ (.A(_03713_),
    .B(_03714_),
    .Y(_03715_));
 sky130_fd_sc_hd__and4_2 _11374_ (.A(_01312_),
    .B(_00544_),
    .C(_01957_),
    .D(_03690_),
    .X(_03716_));
 sky130_fd_sc_hd__and2b_1 _11375_ (.A_N(_03715_),
    .B(_03716_),
    .X(_03717_));
 sky130_fd_sc_hd__o22a_1 _11376_ (.A1(_03695_),
    .A2(_03698_),
    .B1(_03700_),
    .B2(_03692_),
    .X(_03719_));
 sky130_fd_sc_hd__nor2_1 _11377_ (.A(_03701_),
    .B(_03719_),
    .Y(_03720_));
 sky130_fd_sc_hd__nand2_1 _11378_ (.A(_03717_),
    .B(_03720_),
    .Y(_03721_));
 sky130_fd_sc_hd__or3_1 _11379_ (.A(_03711_),
    .B(_03712_),
    .C(_03721_),
    .X(_03722_));
 sky130_fd_sc_hd__and2b_1 _11380_ (.A_N(_03711_),
    .B(_03722_),
    .X(_03723_));
 sky130_fd_sc_hd__a31o_1 _11381_ (.A1(_01312_),
    .A2(_03699_),
    .A3(_03703_),
    .B1(_03702_),
    .X(_03724_));
 sky130_fd_sc_hd__and4_1 _11382_ (.A(_02246_),
    .B(_02249_),
    .C(_03697_),
    .D(_03699_),
    .X(_03725_));
 sky130_fd_sc_hd__a22oi_1 _11383_ (.A1(_02246_),
    .A2(_03697_),
    .B1(_03699_),
    .B2(_02249_),
    .Y(_03726_));
 sky130_fd_sc_hd__nor2_1 _11384_ (.A(_03725_),
    .B(_03726_),
    .Y(_03727_));
 sky130_fd_sc_hd__and2_1 _11385_ (.A(_03724_),
    .B(_03727_),
    .X(_03728_));
 sky130_fd_sc_hd__nor2_1 _11386_ (.A(_03724_),
    .B(_03727_),
    .Y(_03730_));
 sky130_fd_sc_hd__nor2_1 _11387_ (.A(_03728_),
    .B(_03730_),
    .Y(_03731_));
 sky130_fd_sc_hd__xor2_1 _11388_ (.A(_03708_),
    .B(_03731_),
    .X(_03732_));
 sky130_fd_sc_hd__and2b_1 _11389_ (.A_N(_03723_),
    .B(_03732_),
    .X(_03733_));
 sky130_fd_sc_hd__and2b_1 _11390_ (.A_N(_03732_),
    .B(_03723_),
    .X(_03734_));
 sky130_fd_sc_hd__nor2_1 _11391_ (.A(_03733_),
    .B(_03734_),
    .Y(_03735_));
 sky130_fd_sc_hd__and4_1 _11392_ (.A(_00112_),
    .B(_00268_),
    .C(_01179_),
    .D(_01254_),
    .X(_03736_));
 sky130_fd_sc_hd__a22oi_1 _11393_ (.A1(_00113_),
    .A2(_01179_),
    .B1(_01249_),
    .B2(_00114_),
    .Y(_03737_));
 sky130_fd_sc_hd__clkbuf_4 _11394_ (.A(_02119_),
    .X(_03738_));
 sky130_fd_sc_hd__and4bb_1 _11395_ (.A_N(_03736_),
    .B_N(_03737_),
    .C(_06765_),
    .D(_03738_),
    .X(_03739_));
 sky130_fd_sc_hd__and4_1 _11396_ (.A(_00112_),
    .B(_00268_),
    .C(_01254_),
    .D(_02119_),
    .X(_03741_));
 sky130_fd_sc_hd__a22o_1 _11397_ (.A1(_00112_),
    .A2(_01254_),
    .B1(_02119_),
    .B2(_00268_),
    .X(_03742_));
 sky130_fd_sc_hd__and2b_1 _11398_ (.A_N(_03741_),
    .B(_03742_),
    .X(_03743_));
 sky130_fd_sc_hd__clkbuf_4 _11399_ (.A(_02120_),
    .X(_03744_));
 sky130_fd_sc_hd__nand2_1 _11400_ (.A(_00003_),
    .B(_03744_),
    .Y(_03745_));
 sky130_fd_sc_hd__xnor2_1 _11401_ (.A(_03743_),
    .B(_03745_),
    .Y(_03746_));
 sky130_fd_sc_hd__o21ai_2 _11402_ (.A1(_03736_),
    .A2(_03739_),
    .B1(_03746_),
    .Y(_03747_));
 sky130_fd_sc_hd__clkbuf_4 _11403_ (.A(_03744_),
    .X(_03748_));
 sky130_fd_sc_hd__a31o_1 _11404_ (.A1(_00004_),
    .A2(_03748_),
    .A3(_03742_),
    .B1(_03741_),
    .X(_03749_));
 sky130_fd_sc_hd__clkbuf_4 _11405_ (.A(_02119_),
    .X(_03750_));
 sky130_fd_sc_hd__nand4_1 _11406_ (.A(_00257_),
    .B(_00670_),
    .C(_03750_),
    .D(_03748_),
    .Y(_03752_));
 sky130_fd_sc_hd__a22o_1 _11407_ (.A1(_00257_),
    .A2(_03750_),
    .B1(_03748_),
    .B2(_00670_),
    .X(_03753_));
 sky130_fd_sc_hd__and3_1 _11408_ (.A(_03749_),
    .B(_03752_),
    .C(_03753_),
    .X(_03754_));
 sky130_fd_sc_hd__a21oi_1 _11409_ (.A1(_03752_),
    .A2(_03753_),
    .B1(_03749_),
    .Y(_03755_));
 sky130_fd_sc_hd__nor2_1 _11410_ (.A(_03754_),
    .B(_03755_),
    .Y(_03756_));
 sky130_fd_sc_hd__or2b_1 _11411_ (.A(_03747_),
    .B_N(_03756_),
    .X(_03757_));
 sky130_fd_sc_hd__nand4_1 _11412_ (.A(_00114_),
    .B(_06765_),
    .C(_01179_),
    .D(_01254_),
    .Y(_03758_));
 sky130_fd_sc_hd__a22o_1 _11413_ (.A1(_00268_),
    .A2(_01178_),
    .B1(_01248_),
    .B2(_06733_),
    .X(_03759_));
 sky130_fd_sc_hd__nand2_1 _11414_ (.A(_03758_),
    .B(_03759_),
    .Y(_03760_));
 sky130_fd_sc_hd__nand2_1 _11415_ (.A(_06775_),
    .B(_02119_),
    .Y(_03761_));
 sky130_fd_sc_hd__o21ai_1 _11416_ (.A1(_03760_),
    .A2(_03761_),
    .B1(_03758_),
    .Y(_03763_));
 sky130_fd_sc_hd__o2bb2a_1 _11417_ (.A1_N(_00003_),
    .A2_N(_03738_),
    .B1(_03736_),
    .B2(_03737_),
    .X(_03764_));
 sky130_fd_sc_hd__or2_1 _11418_ (.A(_03739_),
    .B(_03764_),
    .X(_03765_));
 sky130_fd_sc_hd__nand2_1 _11419_ (.A(_06775_),
    .B(_03744_),
    .Y(_03766_));
 sky130_fd_sc_hd__xnor2_1 _11420_ (.A(_03763_),
    .B(_03766_),
    .Y(_03767_));
 sky130_fd_sc_hd__and2b_1 _11421_ (.A_N(_03765_),
    .B(_03767_),
    .X(_03768_));
 sky130_fd_sc_hd__a31o_1 _11422_ (.A1(_07004_),
    .A2(_03748_),
    .A3(_03763_),
    .B1(_03768_),
    .X(_03769_));
 sky130_fd_sc_hd__or3_1 _11423_ (.A(_03736_),
    .B(_03739_),
    .C(_03746_),
    .X(_03770_));
 sky130_fd_sc_hd__and2_1 _11424_ (.A(_03747_),
    .B(_03770_),
    .X(_03771_));
 sky130_fd_sc_hd__xnor2_1 _11425_ (.A(_03769_),
    .B(_03771_),
    .Y(_03772_));
 sky130_fd_sc_hd__xor2_1 _11426_ (.A(_03760_),
    .B(_03761_),
    .X(_03774_));
 sky130_fd_sc_hd__and4_1 _11427_ (.A(_00004_),
    .B(_06885_),
    .C(_01180_),
    .D(_01249_),
    .X(_03775_));
 sky130_fd_sc_hd__and2_1 _11428_ (.A(_03774_),
    .B(_03775_),
    .X(_03776_));
 sky130_fd_sc_hd__xnor2_1 _11429_ (.A(_03765_),
    .B(_03767_),
    .Y(_03777_));
 sky130_fd_sc_hd__nand2_1 _11430_ (.A(_03776_),
    .B(_03777_),
    .Y(_03778_));
 sky130_fd_sc_hd__nand2_1 _11431_ (.A(_03769_),
    .B(_03771_),
    .Y(_03779_));
 sky130_fd_sc_hd__o21a_1 _11432_ (.A1(_03772_),
    .A2(_03778_),
    .B1(_03779_),
    .X(_03780_));
 sky130_fd_sc_hd__xnor2_1 _11433_ (.A(_03747_),
    .B(_03756_),
    .Y(_03781_));
 sky130_fd_sc_hd__or2b_1 _11434_ (.A(_03780_),
    .B_N(_03781_),
    .X(_03782_));
 sky130_fd_sc_hd__clkbuf_4 _11435_ (.A(_03748_),
    .X(_03783_));
 sky130_fd_sc_hd__clkbuf_4 _11436_ (.A(_03750_),
    .X(_03785_));
 sky130_fd_sc_hd__nand2_1 _11437_ (.A(_00844_),
    .B(_03785_),
    .Y(_03786_));
 sky130_fd_sc_hd__and3_1 _11438_ (.A(_00843_),
    .B(_03783_),
    .C(_03786_),
    .X(_03787_));
 sky130_fd_sc_hd__xnor2_1 _11439_ (.A(_03754_),
    .B(_03787_),
    .Y(_03788_));
 sky130_fd_sc_hd__a21oi_2 _11440_ (.A1(_03757_),
    .A2(_03782_),
    .B1(_03788_),
    .Y(_03789_));
 sky130_fd_sc_hd__a21bo_1 _11441_ (.A1(_03754_),
    .A2(_03787_),
    .B1_N(_03752_),
    .X(_03790_));
 sky130_fd_sc_hd__a22o_1 _11442_ (.A1(_06964_),
    .A2(_02133_),
    .B1(_02459_),
    .B2(_00121_),
    .X(_03791_));
 sky130_fd_sc_hd__and4_1 _11443_ (.A(_06964_),
    .B(_00121_),
    .C(_02133_),
    .D(_02459_),
    .X(_03792_));
 sky130_fd_sc_hd__a31o_1 _11444_ (.A1(_03554_),
    .A2(_03678_),
    .A3(_03791_),
    .B1(_03792_),
    .X(_03793_));
 sky130_fd_sc_hd__nand4_1 _11445_ (.A(_00262_),
    .B(_00263_),
    .C(_03682_),
    .D(_03679_),
    .Y(_03794_));
 sky130_fd_sc_hd__a22o_1 _11446_ (.A1(_00262_),
    .A2(_03682_),
    .B1(_03678_),
    .B2(_00263_),
    .X(_03796_));
 sky130_fd_sc_hd__and3_1 _11447_ (.A(_03793_),
    .B(_03794_),
    .C(_03796_),
    .X(_03797_));
 sky130_fd_sc_hd__nand2_1 _11448_ (.A(_00263_),
    .B(_03683_),
    .Y(_03798_));
 sky130_fd_sc_hd__and3_1 _11449_ (.A(_00262_),
    .B(_03680_),
    .C(_03798_),
    .X(_03799_));
 sky130_fd_sc_hd__a21bo_1 _11450_ (.A1(_03797_),
    .A2(_03799_),
    .B1_N(_03794_),
    .X(_03800_));
 sky130_fd_sc_hd__and4_1 _11451_ (.A(_06964_),
    .B(_00121_),
    .C(_01953_),
    .D(_02133_),
    .X(_03801_));
 sky130_fd_sc_hd__a22oi_1 _11452_ (.A1(_06964_),
    .A2(_01953_),
    .B1(_02134_),
    .B2(_06966_),
    .Y(_03802_));
 sky130_fd_sc_hd__and4bb_1 _11453_ (.A_N(_03801_),
    .B_N(_03802_),
    .C(_03532_),
    .D(_03681_),
    .X(_03803_));
 sky130_fd_sc_hd__and2b_1 _11454_ (.A_N(_03792_),
    .B(_03791_),
    .X(_03804_));
 sky130_fd_sc_hd__nand2_1 _11455_ (.A(_03543_),
    .B(_02673_),
    .Y(_03805_));
 sky130_fd_sc_hd__xnor2_1 _11456_ (.A(_03804_),
    .B(_03805_),
    .Y(_03807_));
 sky130_fd_sc_hd__o21ai_2 _11457_ (.A1(_03801_),
    .A2(_03803_),
    .B1(_03807_),
    .Y(_03808_));
 sky130_fd_sc_hd__a21oi_1 _11458_ (.A1(_03794_),
    .A2(_03796_),
    .B1(_03793_),
    .Y(_03809_));
 sky130_fd_sc_hd__nor2_1 _11459_ (.A(_03797_),
    .B(_03809_),
    .Y(_03810_));
 sky130_fd_sc_hd__or2b_1 _11460_ (.A(_03808_),
    .B_N(_03810_),
    .X(_03811_));
 sky130_fd_sc_hd__nand4_1 _11461_ (.A(_03532_),
    .B(_00121_),
    .C(_01953_),
    .D(_02134_),
    .Y(_03812_));
 sky130_fd_sc_hd__a22o_1 _11462_ (.A1(_00121_),
    .A2(net21),
    .B1(_02133_),
    .B2(_03521_),
    .X(_03813_));
 sky130_fd_sc_hd__nand2_1 _11463_ (.A(_03812_),
    .B(_03813_),
    .Y(_03814_));
 sky130_fd_sc_hd__nand2_1 _11464_ (.A(_00497_),
    .B(_03681_),
    .Y(_03815_));
 sky130_fd_sc_hd__o21ai_1 _11465_ (.A1(_03814_),
    .A2(_03815_),
    .B1(_03812_),
    .Y(_03816_));
 sky130_fd_sc_hd__o2bb2a_1 _11466_ (.A1_N(_03543_),
    .A2_N(_03681_),
    .B1(_03801_),
    .B2(_03802_),
    .X(_03818_));
 sky130_fd_sc_hd__or2_1 _11467_ (.A(_03803_),
    .B(_03818_),
    .X(_03819_));
 sky130_fd_sc_hd__nand2_1 _11468_ (.A(_00497_),
    .B(_02673_),
    .Y(_03820_));
 sky130_fd_sc_hd__xnor2_1 _11469_ (.A(_03816_),
    .B(_03820_),
    .Y(_03821_));
 sky130_fd_sc_hd__and2b_1 _11470_ (.A_N(_03819_),
    .B(_03821_),
    .X(_03822_));
 sky130_fd_sc_hd__a31o_1 _11471_ (.A1(_00519_),
    .A2(_03679_),
    .A3(_03816_),
    .B1(_03822_),
    .X(_03823_));
 sky130_fd_sc_hd__or3_1 _11472_ (.A(_03801_),
    .B(_03803_),
    .C(_03807_),
    .X(_03824_));
 sky130_fd_sc_hd__and2_1 _11473_ (.A(_03808_),
    .B(_03824_),
    .X(_03825_));
 sky130_fd_sc_hd__xnor2_1 _11474_ (.A(_03823_),
    .B(_03825_),
    .Y(_03826_));
 sky130_fd_sc_hd__xor2_1 _11475_ (.A(_03814_),
    .B(_03815_),
    .X(_03827_));
 sky130_fd_sc_hd__and4_1 _11476_ (.A(_03554_),
    .B(_00508_),
    .C(_01954_),
    .D(_02135_),
    .X(_03829_));
 sky130_fd_sc_hd__and2_1 _11477_ (.A(_03827_),
    .B(_03829_),
    .X(_03830_));
 sky130_fd_sc_hd__xnor2_1 _11478_ (.A(_03819_),
    .B(_03821_),
    .Y(_03831_));
 sky130_fd_sc_hd__nand2_1 _11479_ (.A(_03830_),
    .B(_03831_),
    .Y(_03832_));
 sky130_fd_sc_hd__nand2_1 _11480_ (.A(_03823_),
    .B(_03825_),
    .Y(_03833_));
 sky130_fd_sc_hd__o21a_1 _11481_ (.A1(_03826_),
    .A2(_03832_),
    .B1(_03833_),
    .X(_03834_));
 sky130_fd_sc_hd__xnor2_1 _11482_ (.A(_03808_),
    .B(_03810_),
    .Y(_03835_));
 sky130_fd_sc_hd__or2b_1 _11483_ (.A(_03834_),
    .B_N(_03835_),
    .X(_03836_));
 sky130_fd_sc_hd__xnor2_1 _11484_ (.A(_03797_),
    .B(_03799_),
    .Y(_03837_));
 sky130_fd_sc_hd__a21oi_2 _11485_ (.A1(_03811_),
    .A2(_03836_),
    .B1(_03837_),
    .Y(_03838_));
 sky130_fd_sc_hd__o22ai_4 _11486_ (.A1(_03789_),
    .A2(_03790_),
    .B1(_03800_),
    .B2(_03838_),
    .Y(_03840_));
 sky130_fd_sc_hd__o21ai_1 _11487_ (.A1(_03711_),
    .A2(_03712_),
    .B1(_03721_),
    .Y(_03841_));
 sky130_fd_sc_hd__and2_1 _11488_ (.A(_03722_),
    .B(_03841_),
    .X(_03842_));
 sky130_fd_sc_hd__and2b_1 _11489_ (.A_N(_03840_),
    .B(_03842_),
    .X(_03843_));
 sky130_fd_sc_hd__nand2_1 _11490_ (.A(_03735_),
    .B(_03843_),
    .Y(_03844_));
 sky130_fd_sc_hd__and3_1 _11491_ (.A(_03757_),
    .B(_03782_),
    .C(_03788_),
    .X(_03845_));
 sky130_fd_sc_hd__or2_1 _11492_ (.A(_03789_),
    .B(_03845_),
    .X(_03846_));
 sky130_fd_sc_hd__and3_1 _11493_ (.A(_03811_),
    .B(_03836_),
    .C(_03837_),
    .X(_03847_));
 sky130_fd_sc_hd__or2_1 _11494_ (.A(_03838_),
    .B(_03847_),
    .X(_03848_));
 sky130_fd_sc_hd__nor2_1 _11495_ (.A(_03846_),
    .B(_03848_),
    .Y(_03849_));
 sky130_fd_sc_hd__or4_1 _11496_ (.A(_03789_),
    .B(_03838_),
    .C(_03790_),
    .D(_03800_),
    .X(_03851_));
 sky130_fd_sc_hd__and2_1 _11497_ (.A(_03840_),
    .B(_03851_),
    .X(_03852_));
 sky130_fd_sc_hd__nand2_1 _11498_ (.A(_03849_),
    .B(_03852_),
    .Y(_03853_));
 sky130_fd_sc_hd__or2_1 _11499_ (.A(_03717_),
    .B(_03720_),
    .X(_03854_));
 sky130_fd_sc_hd__nand2_1 _11500_ (.A(_03721_),
    .B(_03854_),
    .Y(_03855_));
 sky130_fd_sc_hd__or2_1 _11501_ (.A(_03849_),
    .B(_03852_),
    .X(_03856_));
 sky130_fd_sc_hd__or2b_1 _11502_ (.A(_03855_),
    .B_N(_03856_),
    .X(_03857_));
 sky130_fd_sc_hd__xor2_1 _11503_ (.A(_03840_),
    .B(_03842_),
    .X(_03858_));
 sky130_fd_sc_hd__a21oi_1 _11504_ (.A1(_03853_),
    .A2(_03857_),
    .B1(_03858_),
    .Y(_03859_));
 sky130_fd_sc_hd__and3_1 _11505_ (.A(_03858_),
    .B(_03853_),
    .C(_03857_),
    .X(_03860_));
 sky130_fd_sc_hd__or2_2 _11506_ (.A(_03859_),
    .B(_03860_),
    .X(_03862_));
 sky130_fd_sc_hd__xnor2_1 _11507_ (.A(_03781_),
    .B(_03780_),
    .Y(_03863_));
 sky130_fd_sc_hd__xnor2_1 _11508_ (.A(_03835_),
    .B(_03834_),
    .Y(_03864_));
 sky130_fd_sc_hd__and2_1 _11509_ (.A(_03863_),
    .B(_03864_),
    .X(_03865_));
 sky130_fd_sc_hd__and2_1 _11510_ (.A(_03846_),
    .B(_03848_),
    .X(_03866_));
 sky130_fd_sc_hd__nor2_1 _11511_ (.A(_03849_),
    .B(_03866_),
    .Y(_03867_));
 sky130_fd_sc_hd__nand2_1 _11512_ (.A(_03865_),
    .B(_03867_),
    .Y(_03868_));
 sky130_fd_sc_hd__xnor2_4 _11513_ (.A(_03715_),
    .B(_03716_),
    .Y(_03869_));
 sky130_fd_sc_hd__or2_1 _11514_ (.A(_03865_),
    .B(_03867_),
    .X(_03870_));
 sky130_fd_sc_hd__nand2_1 _11515_ (.A(_03869_),
    .B(_03870_),
    .Y(_03871_));
 sky130_fd_sc_hd__nand2_1 _11516_ (.A(_03853_),
    .B(_03856_),
    .Y(_03873_));
 sky130_fd_sc_hd__xnor2_1 _11517_ (.A(_03855_),
    .B(_03873_),
    .Y(_03874_));
 sky130_fd_sc_hd__a21o_1 _11518_ (.A1(_03868_),
    .A2(_03871_),
    .B1(_03874_),
    .X(_03875_));
 sky130_fd_sc_hd__nand2_2 _11519_ (.A(_03868_),
    .B(_03870_),
    .Y(_03876_));
 sky130_fd_sc_hd__xor2_4 _11520_ (.A(_03869_),
    .B(_03876_),
    .X(_03877_));
 sky130_fd_sc_hd__xor2_1 _11521_ (.A(_03772_),
    .B(_03778_),
    .X(_03878_));
 sky130_fd_sc_hd__xor2_1 _11522_ (.A(_03826_),
    .B(_03832_),
    .X(_03879_));
 sky130_fd_sc_hd__nand2_1 _11523_ (.A(_03878_),
    .B(_03879_),
    .Y(_03880_));
 sky130_fd_sc_hd__nor2_1 _11524_ (.A(_03863_),
    .B(_03864_),
    .Y(_03881_));
 sky130_fd_sc_hd__or2_1 _11525_ (.A(_03865_),
    .B(_03881_),
    .X(_03882_));
 sky130_fd_sc_hd__nand2_1 _11526_ (.A(_03880_),
    .B(_03882_),
    .Y(_03884_));
 sky130_fd_sc_hd__a22oi_1 _11527_ (.A1(_01312_),
    .A2(_01957_),
    .B1(_03690_),
    .B2(_01155_),
    .Y(_03885_));
 sky130_fd_sc_hd__nor2_1 _11528_ (.A(_03716_),
    .B(_03885_),
    .Y(_03886_));
 sky130_fd_sc_hd__or2_1 _11529_ (.A(_03880_),
    .B(_03882_),
    .X(_03887_));
 sky130_fd_sc_hd__a21bo_2 _11530_ (.A1(_03884_),
    .A2(_03886_),
    .B1_N(_03887_),
    .X(_03888_));
 sky130_fd_sc_hd__xnor2_4 _11531_ (.A(_03877_),
    .B(_03888_),
    .Y(_03889_));
 sky130_fd_sc_hd__nand2_1 _11532_ (.A(_03887_),
    .B(_03884_),
    .Y(_03890_));
 sky130_fd_sc_hd__xor2_2 _11533_ (.A(_03886_),
    .B(_03890_),
    .X(_03891_));
 sky130_fd_sc_hd__or2_1 _11534_ (.A(_03776_),
    .B(_03777_),
    .X(_03892_));
 sky130_fd_sc_hd__and2_1 _11535_ (.A(_03778_),
    .B(_03892_),
    .X(_03893_));
 sky130_fd_sc_hd__and4_1 _11536_ (.A(_06819_),
    .B(_06874_),
    .C(_01177_),
    .D(_01247_),
    .X(_03895_));
 sky130_fd_sc_hd__a22oi_1 _11537_ (.A1(_06873_),
    .A2(_01178_),
    .B1(_01247_),
    .B2(_06874_),
    .Y(_03896_));
 sky130_fd_sc_hd__and4bb_1 _11538_ (.A_N(_03895_),
    .B_N(_03896_),
    .C(_03510_),
    .D(_01564_),
    .X(_03897_));
 sky130_fd_sc_hd__nor2_1 _11539_ (.A(_03895_),
    .B(_03897_),
    .Y(_03898_));
 sky130_fd_sc_hd__and4_1 _11540_ (.A(_06819_),
    .B(_06874_),
    .C(_01247_),
    .D(net19),
    .X(_03899_));
 sky130_fd_sc_hd__a22o_1 _11541_ (.A1(_06873_),
    .A2(_01247_),
    .B1(_01564_),
    .B2(_06874_),
    .X(_03900_));
 sky130_fd_sc_hd__and2b_1 _11542_ (.A_N(_03899_),
    .B(_03900_),
    .X(_03901_));
 sky130_fd_sc_hd__nand2_1 _11543_ (.A(_03521_),
    .B(_01960_),
    .Y(_03902_));
 sky130_fd_sc_hd__xnor2_1 _11544_ (.A(_03901_),
    .B(_03902_),
    .Y(_03903_));
 sky130_fd_sc_hd__or2b_1 _11545_ (.A(_03898_),
    .B_N(_03903_),
    .X(_03904_));
 sky130_fd_sc_hd__a31o_1 _11546_ (.A1(_03532_),
    .A2(_02120_),
    .A3(_03900_),
    .B1(_03899_),
    .X(_03906_));
 sky130_fd_sc_hd__nand4_1 _11547_ (.A(_06965_),
    .B(_06966_),
    .C(_02119_),
    .D(_02120_),
    .Y(_03907_));
 sky130_fd_sc_hd__a22o_1 _11548_ (.A1(_06964_),
    .A2(_02119_),
    .B1(_02120_),
    .B2(_00121_),
    .X(_03908_));
 sky130_fd_sc_hd__and3_1 _11549_ (.A(_03906_),
    .B(_03907_),
    .C(_03908_),
    .X(_03909_));
 sky130_fd_sc_hd__a21oi_1 _11550_ (.A1(_03907_),
    .A2(_03908_),
    .B1(_03906_),
    .Y(_03910_));
 sky130_fd_sc_hd__nor2_1 _11551_ (.A(_03909_),
    .B(_03910_),
    .Y(_03911_));
 sky130_fd_sc_hd__or2b_1 _11552_ (.A(_03904_),
    .B_N(_03911_),
    .X(_03912_));
 sky130_fd_sc_hd__a22o_1 _11553_ (.A1(_06874_),
    .A2(_01177_),
    .B1(_01247_),
    .B2(_03510_),
    .X(_03913_));
 sky130_fd_sc_hd__and3_1 _11554_ (.A(_03510_),
    .B(_06874_),
    .C(_01177_),
    .X(_03914_));
 sky130_fd_sc_hd__a32o_1 _11555_ (.A1(_00486_),
    .A2(_01564_),
    .A3(_03913_),
    .B1(_03914_),
    .B2(_01247_),
    .X(_03915_));
 sky130_fd_sc_hd__and3_1 _11556_ (.A(_00497_),
    .B(_02120_),
    .C(_03915_),
    .X(_03917_));
 sky130_fd_sc_hd__o2bb2a_1 _11557_ (.A1_N(_03521_),
    .A2_N(_02117_),
    .B1(_03895_),
    .B2(_03896_),
    .X(_03918_));
 sky130_fd_sc_hd__or2_1 _11558_ (.A(_03897_),
    .B(_03918_),
    .X(_03919_));
 sky130_fd_sc_hd__nand2_1 _11559_ (.A(_00486_),
    .B(_01960_),
    .Y(_03920_));
 sky130_fd_sc_hd__xnor2_1 _11560_ (.A(_03915_),
    .B(_03920_),
    .Y(_03921_));
 sky130_fd_sc_hd__and2b_1 _11561_ (.A_N(_03919_),
    .B(_03921_),
    .X(_03922_));
 sky130_fd_sc_hd__xnor2_1 _11562_ (.A(_03898_),
    .B(_03903_),
    .Y(_03923_));
 sky130_fd_sc_hd__nor3_1 _11563_ (.A(_03917_),
    .B(_03922_),
    .C(_03923_),
    .Y(_03924_));
 sky130_fd_sc_hd__a21bo_1 _11564_ (.A1(_01247_),
    .A2(_03914_),
    .B1_N(_03913_),
    .X(_03925_));
 sky130_fd_sc_hd__nand2_1 _11565_ (.A(_00486_),
    .B(_02117_),
    .Y(_03926_));
 sky130_fd_sc_hd__xnor2_1 _11566_ (.A(_03925_),
    .B(_03926_),
    .Y(_03928_));
 sky130_fd_sc_hd__and4_1 _11567_ (.A(_03532_),
    .B(_00497_),
    .C(_01179_),
    .D(_01254_),
    .X(_03929_));
 sky130_fd_sc_hd__and2b_1 _11568_ (.A_N(_03928_),
    .B(_03929_),
    .X(_03930_));
 sky130_fd_sc_hd__xnor2_1 _11569_ (.A(_03919_),
    .B(_03921_),
    .Y(_03931_));
 sky130_fd_sc_hd__nand2_1 _11570_ (.A(_03930_),
    .B(_03931_),
    .Y(_03932_));
 sky130_fd_sc_hd__o21a_1 _11571_ (.A1(_03917_),
    .A2(_03922_),
    .B1(_03923_),
    .X(_03933_));
 sky130_fd_sc_hd__o21ba_1 _11572_ (.A1(_03924_),
    .A2(_03932_),
    .B1_N(_03933_),
    .X(_03934_));
 sky130_fd_sc_hd__xnor2_1 _11573_ (.A(_03904_),
    .B(_03911_),
    .Y(_03935_));
 sky130_fd_sc_hd__or2b_1 _11574_ (.A(_03934_),
    .B_N(_03935_),
    .X(_03936_));
 sky130_fd_sc_hd__nand2_1 _11575_ (.A(_00263_),
    .B(_03750_),
    .Y(_03937_));
 sky130_fd_sc_hd__and3_1 _11576_ (.A(_00262_),
    .B(_03748_),
    .C(_03937_),
    .X(_03939_));
 sky130_fd_sc_hd__xnor2_1 _11577_ (.A(_03909_),
    .B(_03939_),
    .Y(_03940_));
 sky130_fd_sc_hd__a21oi_1 _11578_ (.A1(_03912_),
    .A2(_03936_),
    .B1(_03940_),
    .Y(_03941_));
 sky130_fd_sc_hd__a21bo_1 _11579_ (.A1(_03909_),
    .A2(_03939_),
    .B1_N(_03907_),
    .X(_03942_));
 sky130_fd_sc_hd__or3_1 _11580_ (.A(_03893_),
    .B(_03941_),
    .C(_03942_),
    .X(_03943_));
 sky130_fd_sc_hd__o21ai_1 _11581_ (.A1(_03941_),
    .A2(_03942_),
    .B1(_03893_),
    .Y(_03944_));
 sky130_fd_sc_hd__or2_1 _11582_ (.A(_03830_),
    .B(_03831_),
    .X(_03945_));
 sky130_fd_sc_hd__nand2_1 _11583_ (.A(_03832_),
    .B(_03945_),
    .Y(_03946_));
 sky130_fd_sc_hd__nand2_1 _11584_ (.A(_03944_),
    .B(_03946_),
    .Y(_03947_));
 sky130_fd_sc_hd__or2_1 _11585_ (.A(_03878_),
    .B(_03879_),
    .X(_03948_));
 sky130_fd_sc_hd__and2_1 _11586_ (.A(_03880_),
    .B(_03948_),
    .X(_03950_));
 sky130_fd_sc_hd__a21oi_1 _11587_ (.A1(_03943_),
    .A2(_03947_),
    .B1(_03950_),
    .Y(_03951_));
 sky130_fd_sc_hd__and3_1 _11588_ (.A(_03950_),
    .B(_03943_),
    .C(_03947_),
    .X(_03952_));
 sky130_fd_sc_hd__a21oi_1 _11589_ (.A1(_01155_),
    .A2(_01957_),
    .B1(_03952_),
    .Y(_03953_));
 sky130_fd_sc_hd__or2_2 _11590_ (.A(_03951_),
    .B(_03953_),
    .X(_03954_));
 sky130_fd_sc_hd__xor2_1 _11591_ (.A(_03891_),
    .B(_03954_),
    .X(_03955_));
 sky130_fd_sc_hd__inv_2 _11592_ (.A(_03955_),
    .Y(_03956_));
 sky130_fd_sc_hd__nand2_1 _11593_ (.A(_03943_),
    .B(_03944_),
    .Y(_03957_));
 sky130_fd_sc_hd__xor2_1 _11594_ (.A(_03946_),
    .B(_03957_),
    .X(_03958_));
 sky130_fd_sc_hd__nor2_1 _11595_ (.A(_03774_),
    .B(_03775_),
    .Y(_03959_));
 sky130_fd_sc_hd__or2_1 _11596_ (.A(_03776_),
    .B(_03959_),
    .X(_03961_));
 sky130_fd_sc_hd__and3_1 _11597_ (.A(_03940_),
    .B(_03912_),
    .C(_03936_),
    .X(_03962_));
 sky130_fd_sc_hd__or2_1 _11598_ (.A(_03941_),
    .B(_03962_),
    .X(_03963_));
 sky130_fd_sc_hd__nor2_1 _11599_ (.A(_03961_),
    .B(_03963_),
    .Y(_03964_));
 sky130_fd_sc_hd__nor2_1 _11600_ (.A(_03827_),
    .B(_03829_),
    .Y(_03965_));
 sky130_fd_sc_hd__nor2_1 _11601_ (.A(_03830_),
    .B(_03965_),
    .Y(_03966_));
 sky130_fd_sc_hd__nand2_1 _11602_ (.A(_03961_),
    .B(_03963_),
    .Y(_03967_));
 sky130_fd_sc_hd__o21a_1 _11603_ (.A1(_03964_),
    .A2(_03966_),
    .B1(_03967_),
    .X(_03968_));
 sky130_fd_sc_hd__and2_1 _11604_ (.A(_03958_),
    .B(_03968_),
    .X(_03969_));
 sky130_fd_sc_hd__inv_2 _11605_ (.A(_03967_),
    .Y(_03970_));
 sky130_fd_sc_hd__nor2_1 _11606_ (.A(_03970_),
    .B(_03964_),
    .Y(_03972_));
 sky130_fd_sc_hd__xnor2_2 _11607_ (.A(_03966_),
    .B(_03972_),
    .Y(_03973_));
 sky130_fd_sc_hd__inv_2 _11608_ (.A(_03775_),
    .Y(_03974_));
 sky130_fd_sc_hd__a22o_1 _11609_ (.A1(_00654_),
    .A2(_01181_),
    .B1(_01250_),
    .B2(_00543_),
    .X(_03975_));
 sky130_fd_sc_hd__xnor2_1 _11610_ (.A(_03935_),
    .B(_03934_),
    .Y(_03976_));
 sky130_fd_sc_hd__a21o_1 _11611_ (.A1(_03974_),
    .A2(_03975_),
    .B1(_03976_),
    .X(_03977_));
 sky130_fd_sc_hd__a22oi_1 _11612_ (.A1(_03554_),
    .A2(_01956_),
    .B1(_03687_),
    .B2(_00519_),
    .Y(_03978_));
 sky130_fd_sc_hd__nor2_1 _11613_ (.A(_03829_),
    .B(_03978_),
    .Y(_03979_));
 sky130_fd_sc_hd__nand3_1 _11614_ (.A(_03974_),
    .B(_03975_),
    .C(_03976_),
    .Y(_03980_));
 sky130_fd_sc_hd__a21bo_2 _11615_ (.A1(_03977_),
    .A2(_03979_),
    .B1_N(_03980_),
    .X(_03981_));
 sky130_fd_sc_hd__or2b_1 _11616_ (.A(_03973_),
    .B_N(_03981_),
    .X(_03983_));
 sky130_fd_sc_hd__xor2_4 _11617_ (.A(_03981_),
    .B(_03973_),
    .X(_03984_));
 sky130_fd_sc_hd__nor2_1 _11618_ (.A(_03933_),
    .B(_03924_),
    .Y(_03985_));
 sky130_fd_sc_hd__xnor2_1 _11619_ (.A(_03985_),
    .B(_03932_),
    .Y(_03986_));
 sky130_fd_sc_hd__a21o_1 _11620_ (.A1(_00544_),
    .A2(_01182_),
    .B1(_03986_),
    .X(_03987_));
 sky130_fd_sc_hd__and3_1 _11621_ (.A(_00544_),
    .B(_01182_),
    .C(_03986_),
    .X(_03988_));
 sky130_fd_sc_hd__a21o_1 _11622_ (.A1(_00519_),
    .A2(_01957_),
    .B1(_03988_),
    .X(_03989_));
 sky130_fd_sc_hd__nand2_1 _11623_ (.A(_03987_),
    .B(_03989_),
    .Y(_03990_));
 sky130_fd_sc_hd__nand2_1 _11624_ (.A(_03980_),
    .B(_03977_),
    .Y(_03991_));
 sky130_fd_sc_hd__xor2_2 _11625_ (.A(_03979_),
    .B(_03991_),
    .X(_03992_));
 sky130_fd_sc_hd__or3_1 _11626_ (.A(_03984_),
    .B(_03990_),
    .C(_03992_),
    .X(_03994_));
 sky130_fd_sc_hd__nor2_1 _11627_ (.A(_03958_),
    .B(_03968_),
    .Y(_03995_));
 sky130_fd_sc_hd__or2_1 _11628_ (.A(_03969_),
    .B(_03995_),
    .X(_03996_));
 sky130_fd_sc_hd__a21oi_2 _11629_ (.A1(_03983_),
    .A2(_03994_),
    .B1(_03996_),
    .Y(_03997_));
 sky130_fd_sc_hd__o211ai_1 _11630_ (.A1(_03951_),
    .A2(_03952_),
    .B1(_01155_),
    .C1(_01958_),
    .Y(_03998_));
 sky130_fd_sc_hd__a211o_1 _11631_ (.A1(_01155_),
    .A2(_01957_),
    .B1(_03951_),
    .C1(_03952_),
    .X(_03999_));
 sky130_fd_sc_hd__nand2_1 _11632_ (.A(_03998_),
    .B(_03999_),
    .Y(_04000_));
 sky130_fd_sc_hd__o21ai_1 _11633_ (.A1(_03969_),
    .A2(_03997_),
    .B1(_04000_),
    .Y(_04001_));
 sky130_fd_sc_hd__nor2_1 _11634_ (.A(_03956_),
    .B(_04001_),
    .Y(_04002_));
 sky130_fd_sc_hd__o21bai_4 _11635_ (.A1(_03891_),
    .A2(_03954_),
    .B1_N(_04002_),
    .Y(_04003_));
 sky130_fd_sc_hd__and2b_1 _11636_ (.A_N(_03877_),
    .B(_03888_),
    .X(_04005_));
 sky130_fd_sc_hd__a21oi_2 _11637_ (.A1(_03889_),
    .A2(_04003_),
    .B1(_04005_),
    .Y(_04006_));
 sky130_fd_sc_hd__and3_1 _11638_ (.A(_03868_),
    .B(_03874_),
    .C(_03871_),
    .X(_04007_));
 sky130_fd_sc_hd__a21oi_2 _11639_ (.A1(_03875_),
    .A2(_04006_),
    .B1(_04007_),
    .Y(_04008_));
 sky130_fd_sc_hd__and2b_1 _11640_ (.A_N(_03862_),
    .B(_04008_),
    .X(_04009_));
 sky130_fd_sc_hd__or2_1 _11641_ (.A(_03735_),
    .B(_03843_),
    .X(_04010_));
 sky130_fd_sc_hd__and2_1 _11642_ (.A(_03844_),
    .B(_04010_),
    .X(_04011_));
 sky130_fd_sc_hd__o21ai_2 _11643_ (.A1(_03859_),
    .A2(_04009_),
    .B1(_04011_),
    .Y(_04012_));
 sky130_fd_sc_hd__buf_2 _11644_ (.A(_03699_),
    .X(_04013_));
 sky130_fd_sc_hd__buf_2 _11645_ (.A(_03697_),
    .X(_04014_));
 sky130_fd_sc_hd__nand2_1 _11646_ (.A(_02249_),
    .B(_04014_),
    .Y(_04016_));
 sky130_fd_sc_hd__and3_1 _11647_ (.A(_02246_),
    .B(_04013_),
    .C(_04016_),
    .X(_04017_));
 sky130_fd_sc_hd__xor2_1 _11648_ (.A(_03728_),
    .B(_04017_),
    .X(_04018_));
 sky130_fd_sc_hd__a21o_1 _11649_ (.A1(_03708_),
    .A2(_03731_),
    .B1(_03733_),
    .X(_04019_));
 sky130_fd_sc_hd__xnor2_1 _11650_ (.A(_04018_),
    .B(_04019_),
    .Y(_04020_));
 sky130_fd_sc_hd__a21oi_1 _11651_ (.A1(_03844_),
    .A2(_04012_),
    .B1(_04020_),
    .Y(_04021_));
 sky130_fd_sc_hd__and3_1 _11652_ (.A(_04020_),
    .B(_03844_),
    .C(_04012_),
    .X(_04022_));
 sky130_fd_sc_hd__nor2_1 _11653_ (.A(_04021_),
    .B(_04022_),
    .Y(_04023_));
 sky130_fd_sc_hd__inv_2 _11654_ (.A(_04023_),
    .Y(_04024_));
 sky130_fd_sc_hd__xnor2_4 _11655_ (.A(_03889_),
    .B(_04003_),
    .Y(_04025_));
 sky130_fd_sc_hd__or3_1 _11656_ (.A(_04011_),
    .B(_03859_),
    .C(_04009_),
    .X(_04027_));
 sky130_fd_sc_hd__nand2_2 _11657_ (.A(_04012_),
    .B(_04027_),
    .Y(_04028_));
 sky130_fd_sc_hd__xnor2_4 _11658_ (.A(_03862_),
    .B(_04008_),
    .Y(_04029_));
 sky130_fd_sc_hd__and2b_1 _11659_ (.A_N(_04007_),
    .B(_03875_),
    .X(_04030_));
 sky130_fd_sc_hd__xnor2_1 _11660_ (.A(_04006_),
    .B(_04030_),
    .Y(_04031_));
 sky130_fd_sc_hd__nand2_1 _11661_ (.A(_04029_),
    .B(_04031_),
    .Y(_04032_));
 sky130_fd_sc_hd__and3_1 _11662_ (.A(_00258_),
    .B(_06765_),
    .C(_00414_),
    .X(_04033_));
 sky130_fd_sc_hd__a22o_1 _11663_ (.A1(_00258_),
    .A2(_00414_),
    .B1(_00574_),
    .B2(_06765_),
    .X(_04034_));
 sky130_fd_sc_hd__a21bo_1 _11664_ (.A1(_00575_),
    .A2(_04033_),
    .B1_N(_04034_),
    .X(_04035_));
 sky130_fd_sc_hd__nand2_1 _11665_ (.A(_06885_),
    .B(_01601_),
    .Y(_04036_));
 sky130_fd_sc_hd__xnor2_2 _11666_ (.A(_04035_),
    .B(_04036_),
    .Y(_04038_));
 sky130_fd_sc_hd__and4_1 _11667_ (.A(_00004_),
    .B(_06885_),
    .C(_00416_),
    .D(_01288_),
    .X(_04039_));
 sky130_fd_sc_hd__xnor2_2 _11668_ (.A(_04038_),
    .B(_04039_),
    .Y(_04040_));
 sky130_fd_sc_hd__a32o_1 _11669_ (.A1(_06733_),
    .A2(_03773_),
    .A3(_02601_),
    .B1(_02600_),
    .B2(_03696_),
    .X(_04041_));
 sky130_fd_sc_hd__and4_1 _11670_ (.A(_07010_),
    .B(net38),
    .C(_03718_),
    .D(net10),
    .X(_04042_));
 sky130_fd_sc_hd__a22oi_1 _11671_ (.A1(_07010_),
    .A2(_00423_),
    .B1(_03762_),
    .B2(_00101_),
    .Y(_04043_));
 sky130_fd_sc_hd__and4bb_1 _11672_ (.A_N(_04042_),
    .B_N(_04043_),
    .C(_06733_),
    .D(net11),
    .X(_04044_));
 sky130_fd_sc_hd__o2bb2a_1 _11673_ (.A1_N(_06733_),
    .A2_N(_03938_),
    .B1(_04042_),
    .B2(_04043_),
    .X(_04045_));
 sky130_fd_sc_hd__nor2_1 _11674_ (.A(_04044_),
    .B(_04045_),
    .Y(_04046_));
 sky130_fd_sc_hd__nand2_1 _11675_ (.A(_04041_),
    .B(_04046_),
    .Y(_04047_));
 sky130_fd_sc_hd__nand4_1 _11676_ (.A(_00112_),
    .B(_00268_),
    .C(_00755_),
    .D(_01260_),
    .Y(_04049_));
 sky130_fd_sc_hd__a22o_1 _11677_ (.A1(_07010_),
    .A2(_03773_),
    .B1(_01260_),
    .B2(_00268_),
    .X(_04050_));
 sky130_fd_sc_hd__o211a_1 _11678_ (.A1(_04042_),
    .A2(_04044_),
    .B1(_04049_),
    .C1(_04050_),
    .X(_04051_));
 sky130_fd_sc_hd__a211oi_1 _11679_ (.A1(_04049_),
    .A2(_04050_),
    .B1(_04042_),
    .C1(_04044_),
    .Y(_04052_));
 sky130_fd_sc_hd__nor2_1 _11680_ (.A(_04051_),
    .B(_04052_),
    .Y(_04053_));
 sky130_fd_sc_hd__xor2_1 _11681_ (.A(_04047_),
    .B(_04053_),
    .X(_04054_));
 sky130_fd_sc_hd__or2b_1 _11682_ (.A(_02606_),
    .B_N(_02605_),
    .X(_04055_));
 sky130_fd_sc_hd__xnor2_1 _11683_ (.A(_04041_),
    .B(_04046_),
    .Y(_04056_));
 sky130_fd_sc_hd__and3_1 _11684_ (.A(_04055_),
    .B(_02608_),
    .C(_04056_),
    .X(_04057_));
 sky130_fd_sc_hd__a21o_1 _11685_ (.A1(_04055_),
    .A2(_02608_),
    .B1(_04056_),
    .X(_04058_));
 sky130_fd_sc_hd__o31a_1 _11686_ (.A1(_02407_),
    .A2(_02611_),
    .A3(_04057_),
    .B1(_04058_),
    .X(_04060_));
 sky130_fd_sc_hd__xor2_1 _11687_ (.A(_04054_),
    .B(_04060_),
    .X(_04061_));
 sky130_fd_sc_hd__a32o_1 _11688_ (.A1(_03510_),
    .A2(_00734_),
    .A3(_02619_),
    .B1(_02618_),
    .B2(_00413_),
    .X(_04062_));
 sky130_fd_sc_hd__and4_1 _11689_ (.A(_06819_),
    .B(_06821_),
    .C(_00730_),
    .D(net15),
    .X(_04063_));
 sky130_fd_sc_hd__a22oi_1 _11690_ (.A1(_06819_),
    .A2(_00571_),
    .B1(net15),
    .B2(_06874_),
    .Y(_04064_));
 sky130_fd_sc_hd__and4bb_1 _11691_ (.A_N(_04063_),
    .B_N(_04064_),
    .C(_03510_),
    .D(_01211_),
    .X(_04065_));
 sky130_fd_sc_hd__o2bb2a_1 _11692_ (.A1_N(_03510_),
    .A2_N(_01211_),
    .B1(_04063_),
    .B2(_04064_),
    .X(_04066_));
 sky130_fd_sc_hd__nor2_1 _11693_ (.A(_04065_),
    .B(_04066_),
    .Y(_04067_));
 sky130_fd_sc_hd__nand2_1 _11694_ (.A(_04062_),
    .B(_04067_),
    .Y(_04068_));
 sky130_fd_sc_hd__nand4_1 _11695_ (.A(_06964_),
    .B(_06875_),
    .C(_01272_),
    .D(_01211_),
    .Y(_04069_));
 sky130_fd_sc_hd__a22o_1 _11696_ (.A1(_06873_),
    .A2(_01272_),
    .B1(_01211_),
    .B2(_06875_),
    .X(_04071_));
 sky130_fd_sc_hd__o211a_1 _11697_ (.A1(_04063_),
    .A2(_04065_),
    .B1(_04069_),
    .C1(_04071_),
    .X(_04072_));
 sky130_fd_sc_hd__a211oi_1 _11698_ (.A1(_04069_),
    .A2(_04071_),
    .B1(_04063_),
    .C1(_04065_),
    .Y(_04073_));
 sky130_fd_sc_hd__nor2_1 _11699_ (.A(_04072_),
    .B(_04073_),
    .Y(_04074_));
 sky130_fd_sc_hd__xor2_1 _11700_ (.A(_04068_),
    .B(_04074_),
    .X(_04075_));
 sky130_fd_sc_hd__or2b_1 _11701_ (.A(_02625_),
    .B_N(_02624_),
    .X(_04076_));
 sky130_fd_sc_hd__xnor2_1 _11702_ (.A(_04062_),
    .B(_04067_),
    .Y(_04077_));
 sky130_fd_sc_hd__and3_1 _11703_ (.A(_04076_),
    .B(_02627_),
    .C(_04077_),
    .X(_04078_));
 sky130_fd_sc_hd__a21o_1 _11704_ (.A1(_04076_),
    .A2(_02627_),
    .B1(_04077_),
    .X(_04079_));
 sky130_fd_sc_hd__o31a_1 _11705_ (.A1(_02418_),
    .A2(_02629_),
    .A3(_04078_),
    .B1(_04079_),
    .X(_04080_));
 sky130_fd_sc_hd__xor2_1 _11706_ (.A(_04075_),
    .B(_04080_),
    .X(_04082_));
 sky130_fd_sc_hd__nand2_1 _11707_ (.A(_04061_),
    .B(_04082_),
    .Y(_04083_));
 sky130_fd_sc_hd__and3_1 _11708_ (.A(_04041_),
    .B(_04046_),
    .C(_04053_),
    .X(_04084_));
 sky130_fd_sc_hd__nor2_1 _11709_ (.A(_04054_),
    .B(_04060_),
    .Y(_04085_));
 sky130_fd_sc_hd__nand2_1 _11710_ (.A(_00258_),
    .B(_00915_),
    .Y(_04086_));
 sky130_fd_sc_hd__and3_1 _11711_ (.A(_00257_),
    .B(_00916_),
    .C(_04086_),
    .X(_04087_));
 sky130_fd_sc_hd__xor2_1 _11712_ (.A(_04051_),
    .B(_04087_),
    .X(_04088_));
 sky130_fd_sc_hd__o21a_1 _11713_ (.A1(_04084_),
    .A2(_04085_),
    .B1(_04088_),
    .X(_04089_));
 sky130_fd_sc_hd__nor3_1 _11714_ (.A(_04088_),
    .B(_04084_),
    .C(_04085_),
    .Y(_04090_));
 sky130_fd_sc_hd__nor2_1 _11715_ (.A(_04089_),
    .B(_04090_),
    .Y(_04091_));
 sky130_fd_sc_hd__and3_1 _11716_ (.A(_04062_),
    .B(_04067_),
    .C(_04074_),
    .X(_04093_));
 sky130_fd_sc_hd__nor2_1 _11717_ (.A(_04075_),
    .B(_04080_),
    .Y(_04094_));
 sky130_fd_sc_hd__nand2_1 _11718_ (.A(_00263_),
    .B(_01600_),
    .Y(_04095_));
 sky130_fd_sc_hd__and3_1 _11719_ (.A(_00262_),
    .B(_01585_),
    .C(_04095_),
    .X(_04096_));
 sky130_fd_sc_hd__xor2_1 _11720_ (.A(_04072_),
    .B(_04096_),
    .X(_04097_));
 sky130_fd_sc_hd__o21a_1 _11721_ (.A1(_04093_),
    .A2(_04094_),
    .B1(_04097_),
    .X(_04098_));
 sky130_fd_sc_hd__nor3_1 _11722_ (.A(_04097_),
    .B(_04093_),
    .C(_04094_),
    .Y(_04099_));
 sky130_fd_sc_hd__nor2_1 _11723_ (.A(_04098_),
    .B(_04099_),
    .Y(_04100_));
 sky130_fd_sc_hd__xnor2_1 _11724_ (.A(_04091_),
    .B(_04100_),
    .Y(_04101_));
 sky130_fd_sc_hd__nor2_1 _11725_ (.A(_04083_),
    .B(_04101_),
    .Y(_04102_));
 sky130_fd_sc_hd__and2_1 _11726_ (.A(_04083_),
    .B(_04101_),
    .X(_04104_));
 sky130_fd_sc_hd__nor2_1 _11727_ (.A(_04102_),
    .B(_04104_),
    .Y(_04105_));
 sky130_fd_sc_hd__xnor2_2 _11728_ (.A(_04040_),
    .B(_04105_),
    .Y(_04106_));
 sky130_fd_sc_hd__a21oi_1 _11729_ (.A1(_04055_),
    .A2(_02608_),
    .B1(_04056_),
    .Y(_04107_));
 sky130_fd_sc_hd__nor2_1 _11730_ (.A(_04107_),
    .B(_04057_),
    .Y(_04108_));
 sky130_fd_sc_hd__xnor2_1 _11731_ (.A(_02612_),
    .B(_04108_),
    .Y(_04109_));
 sky130_fd_sc_hd__a21oi_1 _11732_ (.A1(_04076_),
    .A2(_02627_),
    .B1(_04077_),
    .Y(_04110_));
 sky130_fd_sc_hd__nor2_1 _11733_ (.A(_04110_),
    .B(_04078_),
    .Y(_04111_));
 sky130_fd_sc_hd__xnor2_1 _11734_ (.A(_02630_),
    .B(_04111_),
    .Y(_04112_));
 sky130_fd_sc_hd__nor2_1 _11735_ (.A(_04109_),
    .B(_04112_),
    .Y(_04113_));
 sky130_fd_sc_hd__or2_1 _11736_ (.A(_04061_),
    .B(_04082_),
    .X(_04115_));
 sky130_fd_sc_hd__and2_1 _11737_ (.A(_04083_),
    .B(_04115_),
    .X(_04116_));
 sky130_fd_sc_hd__or2_1 _11738_ (.A(_04113_),
    .B(_04116_),
    .X(_04117_));
 sky130_fd_sc_hd__a22oi_1 _11739_ (.A1(_00654_),
    .A2(_01188_),
    .B1(_01289_),
    .B2(_00543_),
    .Y(_04118_));
 sky130_fd_sc_hd__nor2_1 _11740_ (.A(_04039_),
    .B(_04118_),
    .Y(_04119_));
 sky130_fd_sc_hd__nand2_1 _11741_ (.A(_04113_),
    .B(_04116_),
    .Y(_04120_));
 sky130_fd_sc_hd__a21bo_1 _11742_ (.A1(_04117_),
    .A2(_04119_),
    .B1_N(_04120_),
    .X(_04121_));
 sky130_fd_sc_hd__xnor2_2 _11743_ (.A(_04106_),
    .B(_04121_),
    .Y(_04122_));
 sky130_fd_sc_hd__nand2_1 _11744_ (.A(_04120_),
    .B(_04117_),
    .Y(_04123_));
 sky130_fd_sc_hd__xor2_1 _11745_ (.A(_04119_),
    .B(_04123_),
    .X(_04124_));
 sky130_fd_sc_hd__nand2_1 _11746_ (.A(_00543_),
    .B(_01188_),
    .Y(_04126_));
 sky130_fd_sc_hd__inv_2 _11747_ (.A(_04126_),
    .Y(_04127_));
 sky130_fd_sc_hd__nand2_1 _11748_ (.A(_02616_),
    .B(_02633_),
    .Y(_04128_));
 sky130_fd_sc_hd__and2_1 _11749_ (.A(_04109_),
    .B(_04112_),
    .X(_04129_));
 sky130_fd_sc_hd__nor2_1 _11750_ (.A(_04113_),
    .B(_04129_),
    .Y(_04130_));
 sky130_fd_sc_hd__and3_1 _11751_ (.A(_02615_),
    .B(_04128_),
    .C(_04130_),
    .X(_04131_));
 sky130_fd_sc_hd__a21oi_1 _11752_ (.A1(_02615_),
    .A2(_04128_),
    .B1(_04130_),
    .Y(_04132_));
 sky130_fd_sc_hd__o21bai_1 _11753_ (.A1(_04127_),
    .A2(_04131_),
    .B1_N(_04132_),
    .Y(_04133_));
 sky130_fd_sc_hd__xor2_1 _11754_ (.A(_04124_),
    .B(_04133_),
    .X(_04134_));
 sky130_fd_sc_hd__or2b_1 _11755_ (.A(_02634_),
    .B_N(_02637_),
    .X(_04135_));
 sky130_fd_sc_hd__a21o_1 _11756_ (.A1(_04135_),
    .A2(_02643_),
    .B1(_02639_),
    .X(_04137_));
 sky130_fd_sc_hd__nor2_1 _11757_ (.A(_04132_),
    .B(_04131_),
    .Y(_04138_));
 sky130_fd_sc_hd__xnor2_2 _11758_ (.A(_04126_),
    .B(_04138_),
    .Y(_04139_));
 sky130_fd_sc_hd__nor2_1 _11759_ (.A(_04124_),
    .B(_04133_),
    .Y(_04140_));
 sky130_fd_sc_hd__a31o_1 _11760_ (.A1(_04134_),
    .A2(_04137_),
    .A3(_04139_),
    .B1(_04140_),
    .X(_04141_));
 sky130_fd_sc_hd__xnor2_2 _11761_ (.A(_04122_),
    .B(_04141_),
    .Y(_04142_));
 sky130_fd_sc_hd__and3_1 _11762_ (.A(_00138_),
    .B(_02018_),
    .C(_01953_),
    .X(_04143_));
 sky130_fd_sc_hd__a22o_1 _11763_ (.A1(_00138_),
    .A2(_01953_),
    .B1(_02134_),
    .B2(_02018_),
    .X(_04144_));
 sky130_fd_sc_hd__a21bo_1 _11764_ (.A1(_02135_),
    .A2(_04143_),
    .B1_N(_04144_),
    .X(_04145_));
 sky130_fd_sc_hd__nand2_1 _11765_ (.A(_02280_),
    .B(_03682_),
    .Y(_04146_));
 sky130_fd_sc_hd__xnor2_2 _11766_ (.A(_04145_),
    .B(_04146_),
    .Y(_04148_));
 sky130_fd_sc_hd__and4_1 _11767_ (.A(_03070_),
    .B(_02335_),
    .C(_01954_),
    .D(_02135_),
    .X(_04149_));
 sky130_fd_sc_hd__xnor2_2 _11768_ (.A(_04148_),
    .B(_04149_),
    .Y(_04150_));
 sky130_fd_sc_hd__a32o_1 _11769_ (.A1(_02007_),
    .A2(_01564_),
    .A3(_02649_),
    .B1(_02648_),
    .B2(_01178_),
    .X(_04151_));
 sky130_fd_sc_hd__and4_1 _11770_ (.A(_05445_),
    .B(_05731_),
    .C(_01246_),
    .D(net19),
    .X(_04152_));
 sky130_fd_sc_hd__a22oi_1 _11771_ (.A1(_05445_),
    .A2(_01246_),
    .B1(net19),
    .B2(_05467_),
    .Y(_04153_));
 sky130_fd_sc_hd__and4bb_1 _11772_ (.A_N(_04152_),
    .B_N(_04153_),
    .C(_01996_),
    .D(net20),
    .X(_04154_));
 sky130_fd_sc_hd__o2bb2a_1 _11773_ (.A1_N(_01996_),
    .A2_N(_01960_),
    .B1(_04152_),
    .B2(_04153_),
    .X(_04155_));
 sky130_fd_sc_hd__nor2_1 _11774_ (.A(_04154_),
    .B(_04155_),
    .Y(_04156_));
 sky130_fd_sc_hd__nand2_1 _11775_ (.A(_04151_),
    .B(_04156_),
    .Y(_04157_));
 sky130_fd_sc_hd__nand4_1 _11776_ (.A(_05456_),
    .B(_05478_),
    .C(_02117_),
    .D(_01960_),
    .Y(_04159_));
 sky130_fd_sc_hd__a22o_1 _11777_ (.A1(_05456_),
    .A2(_02117_),
    .B1(_01960_),
    .B2(_05478_),
    .X(_04160_));
 sky130_fd_sc_hd__o211a_1 _11778_ (.A1(_04152_),
    .A2(_04154_),
    .B1(_04159_),
    .C1(_04160_),
    .X(_04161_));
 sky130_fd_sc_hd__a211oi_1 _11779_ (.A1(_04159_),
    .A2(_04160_),
    .B1(_04152_),
    .C1(_04154_),
    .Y(_04162_));
 sky130_fd_sc_hd__nor2_1 _11780_ (.A(_04161_),
    .B(_04162_),
    .Y(_04163_));
 sky130_fd_sc_hd__xor2_1 _11781_ (.A(_04157_),
    .B(_04163_),
    .X(_04164_));
 sky130_fd_sc_hd__or2b_1 _11782_ (.A(_02655_),
    .B_N(_02654_),
    .X(_04165_));
 sky130_fd_sc_hd__xnor2_1 _11783_ (.A(_04151_),
    .B(_04156_),
    .Y(_04166_));
 sky130_fd_sc_hd__and3_1 _11784_ (.A(_04165_),
    .B(_02657_),
    .C(_04166_),
    .X(_04167_));
 sky130_fd_sc_hd__a21o_1 _11785_ (.A1(_04165_),
    .A2(_02657_),
    .B1(_04166_),
    .X(_04168_));
 sky130_fd_sc_hd__o31a_1 _11786_ (.A1(_02454_),
    .A2(_02659_),
    .A3(_04167_),
    .B1(_04168_),
    .X(_04170_));
 sky130_fd_sc_hd__xor2_1 _11787_ (.A(_04164_),
    .B(_04170_),
    .X(_04171_));
 sky130_fd_sc_hd__a32o_1 _11788_ (.A1(_02127_),
    .A2(net24),
    .A3(_02668_),
    .B1(_02667_),
    .B2(net21),
    .X(_04172_));
 sky130_fd_sc_hd__and4_1 _11789_ (.A(_03850_),
    .B(_01394_),
    .C(net22),
    .D(net24),
    .X(_04173_));
 sky130_fd_sc_hd__a22oi_1 _11790_ (.A1(_01295_),
    .A2(_02133_),
    .B1(net24),
    .B2(_01306_),
    .Y(_04174_));
 sky130_fd_sc_hd__and4bb_1 _11791_ (.A_N(_04173_),
    .B_N(_04174_),
    .C(_01744_),
    .D(net25),
    .X(_04175_));
 sky130_fd_sc_hd__o2bb2a_1 _11792_ (.A1_N(_02127_),
    .A2_N(net25),
    .B1(_04173_),
    .B2(_04174_),
    .X(_04176_));
 sky130_fd_sc_hd__nor2_1 _11793_ (.A(_04175_),
    .B(_04176_),
    .Y(_04177_));
 sky130_fd_sc_hd__nand2_1 _11794_ (.A(_04172_),
    .B(_04177_),
    .Y(_04178_));
 sky130_fd_sc_hd__nand4_1 _11795_ (.A(_01361_),
    .B(_00159_),
    .C(_02459_),
    .D(_02673_),
    .Y(_04179_));
 sky130_fd_sc_hd__a22o_1 _11796_ (.A1(_01361_),
    .A2(_02459_),
    .B1(_02673_),
    .B2(_01405_),
    .X(_04181_));
 sky130_fd_sc_hd__o211a_1 _11797_ (.A1(_04173_),
    .A2(_04175_),
    .B1(_04179_),
    .C1(_04181_),
    .X(_04182_));
 sky130_fd_sc_hd__a211oi_1 _11798_ (.A1(_04179_),
    .A2(_04181_),
    .B1(_04173_),
    .C1(_04175_),
    .Y(_04183_));
 sky130_fd_sc_hd__nor2_1 _11799_ (.A(_04182_),
    .B(_04183_),
    .Y(_04184_));
 sky130_fd_sc_hd__xor2_1 _11800_ (.A(_04178_),
    .B(_04184_),
    .X(_04185_));
 sky130_fd_sc_hd__or2b_1 _11801_ (.A(_02674_),
    .B_N(_02672_),
    .X(_04186_));
 sky130_fd_sc_hd__xnor2_1 _11802_ (.A(_04172_),
    .B(_04177_),
    .Y(_04187_));
 sky130_fd_sc_hd__and3_1 _11803_ (.A(_04186_),
    .B(_02677_),
    .C(_04187_),
    .X(_04188_));
 sky130_fd_sc_hd__a21o_1 _11804_ (.A1(_04186_),
    .A2(_02677_),
    .B1(_04187_),
    .X(_04189_));
 sky130_fd_sc_hd__o31a_1 _11805_ (.A1(_02466_),
    .A2(_02679_),
    .A3(_04188_),
    .B1(_04189_),
    .X(_04190_));
 sky130_fd_sc_hd__xor2_1 _11806_ (.A(_04185_),
    .B(_04190_),
    .X(_04192_));
 sky130_fd_sc_hd__nand2_1 _11807_ (.A(_04171_),
    .B(_04192_),
    .Y(_04193_));
 sky130_fd_sc_hd__and3_1 _11808_ (.A(_04151_),
    .B(_04156_),
    .C(_04163_),
    .X(_04194_));
 sky130_fd_sc_hd__nor2_1 _11809_ (.A(_04164_),
    .B(_04170_),
    .Y(_04195_));
 sky130_fd_sc_hd__nand2_1 _11810_ (.A(_06439_),
    .B(_03750_),
    .Y(_04196_));
 sky130_fd_sc_hd__and3_1 _11811_ (.A(_06428_),
    .B(_03748_),
    .C(_04196_),
    .X(_04197_));
 sky130_fd_sc_hd__xor2_1 _11812_ (.A(_04161_),
    .B(_04197_),
    .X(_04198_));
 sky130_fd_sc_hd__o21a_1 _11813_ (.A1(_04194_),
    .A2(_04195_),
    .B1(_04198_),
    .X(_04199_));
 sky130_fd_sc_hd__nor3_1 _11814_ (.A(_04198_),
    .B(_04194_),
    .C(_04195_),
    .Y(_04200_));
 sky130_fd_sc_hd__nor2_1 _11815_ (.A(_04199_),
    .B(_04200_),
    .Y(_04201_));
 sky130_fd_sc_hd__and3_1 _11816_ (.A(_04172_),
    .B(_04177_),
    .C(_04184_),
    .X(_04203_));
 sky130_fd_sc_hd__nor2_1 _11817_ (.A(_04185_),
    .B(_04190_),
    .Y(_04204_));
 sky130_fd_sc_hd__nand2_1 _11818_ (.A(_00159_),
    .B(_03682_),
    .Y(_04205_));
 sky130_fd_sc_hd__and3_1 _11819_ (.A(_00157_),
    .B(_03678_),
    .C(_04205_),
    .X(_04206_));
 sky130_fd_sc_hd__xor2_1 _11820_ (.A(_04182_),
    .B(_04206_),
    .X(_04207_));
 sky130_fd_sc_hd__o21a_1 _11821_ (.A1(_04203_),
    .A2(_04204_),
    .B1(_04207_),
    .X(_04208_));
 sky130_fd_sc_hd__nor3_1 _11822_ (.A(_04207_),
    .B(_04203_),
    .C(_04204_),
    .Y(_04209_));
 sky130_fd_sc_hd__nor2_1 _11823_ (.A(_04208_),
    .B(_04209_),
    .Y(_04210_));
 sky130_fd_sc_hd__xnor2_1 _11824_ (.A(_04201_),
    .B(_04210_),
    .Y(_04211_));
 sky130_fd_sc_hd__nor2_1 _11825_ (.A(_04193_),
    .B(_04211_),
    .Y(_04212_));
 sky130_fd_sc_hd__and2_1 _11826_ (.A(_04193_),
    .B(_04211_),
    .X(_04214_));
 sky130_fd_sc_hd__nor2_1 _11827_ (.A(_04212_),
    .B(_04214_),
    .Y(_04215_));
 sky130_fd_sc_hd__xnor2_2 _11828_ (.A(_04150_),
    .B(_04215_),
    .Y(_04216_));
 sky130_fd_sc_hd__a21oi_1 _11829_ (.A1(_04165_),
    .A2(_02657_),
    .B1(_04166_),
    .Y(_04217_));
 sky130_fd_sc_hd__nor2_1 _11830_ (.A(_04217_),
    .B(_04167_),
    .Y(_04218_));
 sky130_fd_sc_hd__xnor2_1 _11831_ (.A(_02660_),
    .B(_04218_),
    .Y(_04219_));
 sky130_fd_sc_hd__a21oi_1 _11832_ (.A1(_04186_),
    .A2(_02677_),
    .B1(_04187_),
    .Y(_04220_));
 sky130_fd_sc_hd__nor2_1 _11833_ (.A(_04220_),
    .B(_04188_),
    .Y(_04221_));
 sky130_fd_sc_hd__xnor2_1 _11834_ (.A(_02680_),
    .B(_04221_),
    .Y(_04222_));
 sky130_fd_sc_hd__nor2_1 _11835_ (.A(_04219_),
    .B(_04222_),
    .Y(_04223_));
 sky130_fd_sc_hd__or2_1 _11836_ (.A(_04171_),
    .B(_04192_),
    .X(_04225_));
 sky130_fd_sc_hd__and2_1 _11837_ (.A(_04193_),
    .B(_04225_),
    .X(_04226_));
 sky130_fd_sc_hd__or2_1 _11838_ (.A(_04223_),
    .B(_04226_),
    .X(_04227_));
 sky130_fd_sc_hd__a22oi_1 _11839_ (.A1(_03070_),
    .A2(_01955_),
    .B1(_03686_),
    .B2(_02456_),
    .Y(_04228_));
 sky130_fd_sc_hd__nor2_1 _11840_ (.A(_04149_),
    .B(_04228_),
    .Y(_04229_));
 sky130_fd_sc_hd__nand2_1 _11841_ (.A(_04223_),
    .B(_04226_),
    .Y(_04230_));
 sky130_fd_sc_hd__a21bo_1 _11842_ (.A1(_04227_),
    .A2(_04229_),
    .B1_N(_04230_),
    .X(_04231_));
 sky130_fd_sc_hd__xnor2_2 _11843_ (.A(_04216_),
    .B(_04231_),
    .Y(_04232_));
 sky130_fd_sc_hd__nand2_1 _11844_ (.A(_04230_),
    .B(_04227_),
    .Y(_04233_));
 sky130_fd_sc_hd__xor2_1 _11845_ (.A(_04229_),
    .B(_04233_),
    .X(_04234_));
 sky130_fd_sc_hd__nand2_2 _11846_ (.A(_02456_),
    .B(_01955_),
    .Y(_04236_));
 sky130_fd_sc_hd__inv_2 _11847_ (.A(_04236_),
    .Y(_04237_));
 sky130_fd_sc_hd__nand2_1 _11848_ (.A(_02665_),
    .B(_02682_),
    .Y(_04238_));
 sky130_fd_sc_hd__and2_1 _11849_ (.A(_04219_),
    .B(_04222_),
    .X(_04239_));
 sky130_fd_sc_hd__nor2_1 _11850_ (.A(_04223_),
    .B(_04239_),
    .Y(_04240_));
 sky130_fd_sc_hd__and3_1 _11851_ (.A(_02663_),
    .B(_04238_),
    .C(_04240_),
    .X(_04241_));
 sky130_fd_sc_hd__a21oi_1 _11852_ (.A1(_02663_),
    .A2(_04238_),
    .B1(_04240_),
    .Y(_04242_));
 sky130_fd_sc_hd__o21bai_1 _11853_ (.A1(_04237_),
    .A2(_04241_),
    .B1_N(_04242_),
    .Y(_04243_));
 sky130_fd_sc_hd__xor2_1 _11854_ (.A(_04234_),
    .B(_04243_),
    .X(_04244_));
 sky130_fd_sc_hd__or2b_1 _11855_ (.A(_02683_),
    .B_N(_02687_),
    .X(_04245_));
 sky130_fd_sc_hd__a21o_1 _11856_ (.A1(_04245_),
    .A2(_02692_),
    .B1(_02689_),
    .X(_04247_));
 sky130_fd_sc_hd__nor2_1 _11857_ (.A(_04242_),
    .B(_04241_),
    .Y(_04248_));
 sky130_fd_sc_hd__xnor2_2 _11858_ (.A(_04236_),
    .B(_04248_),
    .Y(_04249_));
 sky130_fd_sc_hd__nor2_1 _11859_ (.A(_04234_),
    .B(_04243_),
    .Y(_04250_));
 sky130_fd_sc_hd__a31o_1 _11860_ (.A1(_04244_),
    .A2(_04247_),
    .A3(_04249_),
    .B1(_04250_),
    .X(_04251_));
 sky130_fd_sc_hd__xnor2_2 _11861_ (.A(_04232_),
    .B(_04251_),
    .Y(_04252_));
 sky130_fd_sc_hd__nor2_1 _11862_ (.A(_04142_),
    .B(_04252_),
    .Y(_04253_));
 sky130_fd_sc_hd__and2b_1 _11863_ (.A_N(_04106_),
    .B(_04121_),
    .X(_04254_));
 sky130_fd_sc_hd__a21o_1 _11864_ (.A1(_04122_),
    .A2(_04141_),
    .B1(_04254_),
    .X(_04255_));
 sky130_fd_sc_hd__and2b_1 _11865_ (.A_N(_04038_),
    .B(_04039_),
    .X(_04256_));
 sky130_fd_sc_hd__and4_1 _11866_ (.A(_00113_),
    .B(_00258_),
    .C(_00415_),
    .D(_00574_),
    .X(_04258_));
 sky130_fd_sc_hd__a22oi_1 _11867_ (.A1(_00113_),
    .A2(_00415_),
    .B1(_00575_),
    .B2(_00258_),
    .Y(_04259_));
 sky130_fd_sc_hd__and4bb_1 _11868_ (.A_N(_04258_),
    .B_N(_04259_),
    .C(_00003_),
    .D(_01600_),
    .X(_04260_));
 sky130_fd_sc_hd__a32o_1 _11869_ (.A1(_06775_),
    .A2(_01600_),
    .A3(_04034_),
    .B1(_04033_),
    .B2(_00575_),
    .X(_04261_));
 sky130_fd_sc_hd__and3_1 _11870_ (.A(_06885_),
    .B(_01780_),
    .C(_04261_),
    .X(_04262_));
 sky130_fd_sc_hd__o2bb2a_1 _11871_ (.A1_N(_00004_),
    .A2_N(_01601_),
    .B1(_04258_),
    .B2(_04259_),
    .X(_04263_));
 sky130_fd_sc_hd__a21oi_1 _11872_ (.A1(_07004_),
    .A2(_01780_),
    .B1(_04261_),
    .Y(_04264_));
 sky130_fd_sc_hd__nor4_1 _11873_ (.A(_04260_),
    .B(_04262_),
    .C(_04263_),
    .D(_04264_),
    .Y(_04265_));
 sky130_fd_sc_hd__o22a_1 _11874_ (.A1(_04260_),
    .A2(_04263_),
    .B1(_04264_),
    .B2(_04262_),
    .X(_04266_));
 sky130_fd_sc_hd__nor2_1 _11875_ (.A(net146),
    .B(_04266_),
    .Y(_04267_));
 sky130_fd_sc_hd__nand2_1 _11876_ (.A(_04256_),
    .B(_04267_),
    .Y(_04269_));
 sky130_fd_sc_hd__or2_1 _11877_ (.A(_04256_),
    .B(_04267_),
    .X(_04270_));
 sky130_fd_sc_hd__and2_1 _11878_ (.A(_04269_),
    .B(_04270_),
    .X(_04271_));
 sky130_fd_sc_hd__nand2_1 _11879_ (.A(_04091_),
    .B(_04100_),
    .Y(_04272_));
 sky130_fd_sc_hd__and4_1 _11880_ (.A(_00257_),
    .B(_00670_),
    .C(_00915_),
    .D(_00916_),
    .X(_04273_));
 sky130_fd_sc_hd__a211o_1 _11881_ (.A1(_04051_),
    .A2(_04087_),
    .B1(_04089_),
    .C1(_04273_),
    .X(_04274_));
 sky130_fd_sc_hd__and4_1 _11882_ (.A(_00262_),
    .B(_00263_),
    .C(_02090_),
    .D(_01780_),
    .X(_04275_));
 sky130_fd_sc_hd__a211o_1 _11883_ (.A1(_04072_),
    .A2(_04096_),
    .B1(_04098_),
    .C1(_04275_),
    .X(_04276_));
 sky130_fd_sc_hd__xnor2_1 _11884_ (.A(_04274_),
    .B(_04276_),
    .Y(_04277_));
 sky130_fd_sc_hd__nor2_1 _11885_ (.A(_04272_),
    .B(_04277_),
    .Y(_04278_));
 sky130_fd_sc_hd__nand2_1 _11886_ (.A(_04272_),
    .B(_04277_),
    .Y(_04280_));
 sky130_fd_sc_hd__or2b_1 _11887_ (.A(_04278_),
    .B_N(_04280_),
    .X(_04281_));
 sky130_fd_sc_hd__xnor2_1 _11888_ (.A(_04271_),
    .B(_04281_),
    .Y(_04282_));
 sky130_fd_sc_hd__and2b_1 _11889_ (.A_N(_04104_),
    .B(_04040_),
    .X(_04283_));
 sky130_fd_sc_hd__nor3_1 _11890_ (.A(_04282_),
    .B(_04102_),
    .C(_04283_),
    .Y(_04284_));
 sky130_fd_sc_hd__o21a_1 _11891_ (.A1(_04102_),
    .A2(_04283_),
    .B1(_04282_),
    .X(_04285_));
 sky130_fd_sc_hd__nor2_1 _11892_ (.A(_04284_),
    .B(_04285_),
    .Y(_04286_));
 sky130_fd_sc_hd__xnor2_2 _11893_ (.A(_04255_),
    .B(_04286_),
    .Y(_04287_));
 sky130_fd_sc_hd__and2b_1 _11894_ (.A_N(_04216_),
    .B(_04231_),
    .X(_04288_));
 sky130_fd_sc_hd__a21oi_1 _11895_ (.A1(_04232_),
    .A2(_04251_),
    .B1(_04288_),
    .Y(_04289_));
 sky130_fd_sc_hd__and2b_1 _11896_ (.A_N(_04148_),
    .B(_04149_),
    .X(_04291_));
 sky130_fd_sc_hd__and4_1 _11897_ (.A(_06417_),
    .B(_06439_),
    .C(_01954_),
    .D(_02135_),
    .X(_04292_));
 sky130_fd_sc_hd__a22oi_1 _11898_ (.A1(_06428_),
    .A2(_01954_),
    .B1(_02135_),
    .B2(_06439_),
    .Y(_04293_));
 sky130_fd_sc_hd__and4bb_1 _11899_ (.A_N(_04292_),
    .B_N(_04293_),
    .C(_03059_),
    .D(_03682_),
    .X(_04294_));
 sky130_fd_sc_hd__a32o_1 _11900_ (.A1(_02040_),
    .A2(_03681_),
    .A3(_04144_),
    .B1(_04143_),
    .B2(_02135_),
    .X(_04295_));
 sky130_fd_sc_hd__and3_1 _11901_ (.A(_02280_),
    .B(_03678_),
    .C(_04295_),
    .X(_04296_));
 sky130_fd_sc_hd__o2bb2a_1 _11902_ (.A1_N(_03070_),
    .A2_N(_03682_),
    .B1(_04292_),
    .B2(_04293_),
    .X(_04297_));
 sky130_fd_sc_hd__a21oi_1 _11903_ (.A1(_02335_),
    .A2(_03678_),
    .B1(_04295_),
    .Y(_04298_));
 sky130_fd_sc_hd__nor4_1 _11904_ (.A(_04294_),
    .B(_04296_),
    .C(_04297_),
    .D(_04298_),
    .Y(_04299_));
 sky130_fd_sc_hd__o22a_1 _11905_ (.A1(_04294_),
    .A2(_04297_),
    .B1(_04298_),
    .B2(_04296_),
    .X(_04300_));
 sky130_fd_sc_hd__nor2_1 _11906_ (.A(_04299_),
    .B(_04300_),
    .Y(_04302_));
 sky130_fd_sc_hd__nand2_1 _11907_ (.A(_04291_),
    .B(_04302_),
    .Y(_04303_));
 sky130_fd_sc_hd__or2_1 _11908_ (.A(_04291_),
    .B(_04302_),
    .X(_04304_));
 sky130_fd_sc_hd__and2_1 _11909_ (.A(_04303_),
    .B(_04304_),
    .X(_04305_));
 sky130_fd_sc_hd__nand2_1 _11910_ (.A(_04201_),
    .B(_04210_),
    .Y(_04306_));
 sky130_fd_sc_hd__and4_1 _11911_ (.A(_06626_),
    .B(_06450_),
    .C(_03750_),
    .D(_03783_),
    .X(_04307_));
 sky130_fd_sc_hd__a211o_1 _11912_ (.A1(_04161_),
    .A2(_04197_),
    .B1(_04199_),
    .C1(_04307_),
    .X(_04308_));
 sky130_fd_sc_hd__and4_1 _11913_ (.A(_00157_),
    .B(_00159_),
    .C(_03683_),
    .D(_03679_),
    .X(_04309_));
 sky130_fd_sc_hd__a211o_1 _11914_ (.A1(_04182_),
    .A2(_04206_),
    .B1(_04208_),
    .C1(_04309_),
    .X(_04310_));
 sky130_fd_sc_hd__xnor2_1 _11915_ (.A(_04308_),
    .B(_04310_),
    .Y(_04311_));
 sky130_fd_sc_hd__nor2_1 _11916_ (.A(_04306_),
    .B(_04311_),
    .Y(_04313_));
 sky130_fd_sc_hd__nand2_1 _11917_ (.A(_04306_),
    .B(_04311_),
    .Y(_04314_));
 sky130_fd_sc_hd__or2b_1 _11918_ (.A(_04313_),
    .B_N(_04314_),
    .X(_04315_));
 sky130_fd_sc_hd__xnor2_1 _11919_ (.A(_04305_),
    .B(_04315_),
    .Y(_04316_));
 sky130_fd_sc_hd__and2b_1 _11920_ (.A_N(_04214_),
    .B(_04150_),
    .X(_04317_));
 sky130_fd_sc_hd__nor3_1 _11921_ (.A(_04316_),
    .B(_04212_),
    .C(_04317_),
    .Y(_04318_));
 sky130_fd_sc_hd__o21a_1 _11922_ (.A1(_04212_),
    .A2(_04317_),
    .B1(_04316_),
    .X(_04319_));
 sky130_fd_sc_hd__nor2_1 _11923_ (.A(_04318_),
    .B(_04319_),
    .Y(_04320_));
 sky130_fd_sc_hd__xnor2_2 _11924_ (.A(_04289_),
    .B(_04320_),
    .Y(_04321_));
 sky130_fd_sc_hd__xnor2_2 _11925_ (.A(_04287_),
    .B(_04321_),
    .Y(_04322_));
 sky130_fd_sc_hd__nand2_1 _11926_ (.A(_04253_),
    .B(_04322_),
    .Y(_04324_));
 sky130_fd_sc_hd__or2_1 _11927_ (.A(_03930_),
    .B(_03931_),
    .X(_04325_));
 sky130_fd_sc_hd__nand2_1 _11928_ (.A(_03932_),
    .B(_04325_),
    .Y(_04326_));
 sky130_fd_sc_hd__nor2_1 _11929_ (.A(_04253_),
    .B(_04322_),
    .Y(_04327_));
 sky130_fd_sc_hd__a21o_1 _11930_ (.A1(_04324_),
    .A2(_04326_),
    .B1(_04327_),
    .X(_04328_));
 sky130_fd_sc_hd__and4_1 _11931_ (.A(_00113_),
    .B(_00114_),
    .C(_00572_),
    .D(_01272_),
    .X(_04329_));
 sky130_fd_sc_hd__nand2_1 _11932_ (.A(_00114_),
    .B(_01272_),
    .Y(_04330_));
 sky130_fd_sc_hd__a21boi_1 _11933_ (.A1(_00113_),
    .A2(_00574_),
    .B1_N(_04330_),
    .Y(_04331_));
 sky130_fd_sc_hd__nor2_1 _11934_ (.A(_04329_),
    .B(_04331_),
    .Y(_04332_));
 sky130_fd_sc_hd__and3_1 _11935_ (.A(_00003_),
    .B(_01585_),
    .C(_04332_),
    .X(_04333_));
 sky130_fd_sc_hd__a21oi_1 _11936_ (.A1(_00004_),
    .A2(_01585_),
    .B1(_04332_),
    .Y(_04335_));
 sky130_fd_sc_hd__nor2_1 _11937_ (.A(_04333_),
    .B(_04335_),
    .Y(_04336_));
 sky130_fd_sc_hd__o21a_1 _11938_ (.A1(_04258_),
    .A2(_04260_),
    .B1(_04336_),
    .X(_04337_));
 sky130_fd_sc_hd__nor3_1 _11939_ (.A(_04258_),
    .B(_04260_),
    .C(_04336_),
    .Y(_04338_));
 sky130_fd_sc_hd__nor2_1 _11940_ (.A(_04337_),
    .B(_04338_),
    .Y(_04339_));
 sky130_fd_sc_hd__o21a_1 _11941_ (.A1(_04262_),
    .A2(net146),
    .B1(_04339_),
    .X(_04340_));
 sky130_fd_sc_hd__nor3_1 _11942_ (.A(_04262_),
    .B(_04265_),
    .C(_04339_),
    .Y(_04341_));
 sky130_fd_sc_hd__or3_1 _11943_ (.A(_04340_),
    .B(_04269_),
    .C(_04341_),
    .X(_04342_));
 sky130_fd_sc_hd__o21ai_1 _11944_ (.A1(_04340_),
    .A2(_04341_),
    .B1(_04269_),
    .Y(_04343_));
 sky130_fd_sc_hd__and2_1 _11945_ (.A(_04342_),
    .B(_04343_),
    .X(_04344_));
 sky130_fd_sc_hd__and3_1 _11946_ (.A(_04274_),
    .B(_04276_),
    .C(_04344_),
    .X(_04346_));
 sky130_fd_sc_hd__and2_1 _11947_ (.A(_04274_),
    .B(_04276_),
    .X(_04347_));
 sky130_fd_sc_hd__nor2_1 _11948_ (.A(_04347_),
    .B(_04344_),
    .Y(_04348_));
 sky130_fd_sc_hd__or2_1 _11949_ (.A(_04346_),
    .B(_04348_),
    .X(_04349_));
 sky130_fd_sc_hd__a21oi_1 _11950_ (.A1(_04271_),
    .A2(_04280_),
    .B1(_04278_),
    .Y(_04350_));
 sky130_fd_sc_hd__nor2_1 _11951_ (.A(_04349_),
    .B(_04350_),
    .Y(_04351_));
 sky130_fd_sc_hd__and2_1 _11952_ (.A(_04349_),
    .B(_04350_),
    .X(_04352_));
 sky130_fd_sc_hd__nor2_1 _11953_ (.A(_04351_),
    .B(_04352_),
    .Y(_04353_));
 sky130_fd_sc_hd__or3_2 _11954_ (.A(_04282_),
    .B(_04102_),
    .C(_04283_),
    .X(_04354_));
 sky130_fd_sc_hd__a211o_1 _11955_ (.A1(_04122_),
    .A2(_04141_),
    .B1(_04285_),
    .C1(_04254_),
    .X(_04355_));
 sky130_fd_sc_hd__nand3_2 _11956_ (.A(_04353_),
    .B(_04354_),
    .C(_04355_),
    .Y(_04357_));
 sky130_fd_sc_hd__and4_1 _11957_ (.A(_06417_),
    .B(_00138_),
    .C(_02134_),
    .D(_03681_),
    .X(_04358_));
 sky130_fd_sc_hd__nand2_1 _11958_ (.A(_00138_),
    .B(_02459_),
    .Y(_04359_));
 sky130_fd_sc_hd__a21boi_1 _11959_ (.A1(_06417_),
    .A2(_02134_),
    .B1_N(_04359_),
    .Y(_04360_));
 sky130_fd_sc_hd__nor2_1 _11960_ (.A(_04358_),
    .B(_04360_),
    .Y(_04361_));
 sky130_fd_sc_hd__and3_1 _11961_ (.A(_03059_),
    .B(_03678_),
    .C(_04361_),
    .X(_04362_));
 sky130_fd_sc_hd__a21oi_1 _11962_ (.A1(_03059_),
    .A2(_03678_),
    .B1(_04361_),
    .Y(_04363_));
 sky130_fd_sc_hd__nor2_1 _11963_ (.A(_04362_),
    .B(_04363_),
    .Y(_04364_));
 sky130_fd_sc_hd__o21a_1 _11964_ (.A1(_04292_),
    .A2(_04294_),
    .B1(_04364_),
    .X(_04365_));
 sky130_fd_sc_hd__nor3_1 _11965_ (.A(_04292_),
    .B(_04294_),
    .C(_04364_),
    .Y(_04366_));
 sky130_fd_sc_hd__nor2_1 _11966_ (.A(_04365_),
    .B(_04366_),
    .Y(_04368_));
 sky130_fd_sc_hd__o21a_1 _11967_ (.A1(_04296_),
    .A2(net144),
    .B1(_04368_),
    .X(_04369_));
 sky130_fd_sc_hd__nor3_1 _11968_ (.A(_04296_),
    .B(net144),
    .C(_04368_),
    .Y(_04370_));
 sky130_fd_sc_hd__or3_1 _11969_ (.A(_04369_),
    .B(_04303_),
    .C(_04370_),
    .X(_04371_));
 sky130_fd_sc_hd__o21ai_1 _11970_ (.A1(_04369_),
    .A2(_04370_),
    .B1(_04303_),
    .Y(_04372_));
 sky130_fd_sc_hd__and2_1 _11971_ (.A(_04371_),
    .B(_04372_),
    .X(_04373_));
 sky130_fd_sc_hd__and3_1 _11972_ (.A(_04308_),
    .B(_04310_),
    .C(_04373_),
    .X(_04374_));
 sky130_fd_sc_hd__and2_1 _11973_ (.A(_04308_),
    .B(_04310_),
    .X(_04375_));
 sky130_fd_sc_hd__nor2_1 _11974_ (.A(_04375_),
    .B(_04373_),
    .Y(_04376_));
 sky130_fd_sc_hd__or2_1 _11975_ (.A(_04374_),
    .B(_04376_),
    .X(_04377_));
 sky130_fd_sc_hd__a21oi_1 _11976_ (.A1(_04305_),
    .A2(_04314_),
    .B1(_04313_),
    .Y(_04379_));
 sky130_fd_sc_hd__nor2_1 _11977_ (.A(_04377_),
    .B(_04379_),
    .Y(_04380_));
 sky130_fd_sc_hd__and2_1 _11978_ (.A(_04377_),
    .B(_04379_),
    .X(_04381_));
 sky130_fd_sc_hd__nor2_1 _11979_ (.A(_04380_),
    .B(_04381_),
    .Y(_04382_));
 sky130_fd_sc_hd__or3_2 _11980_ (.A(_04316_),
    .B(_04212_),
    .C(_04317_),
    .X(_04383_));
 sky130_fd_sc_hd__a211o_1 _11981_ (.A1(_04232_),
    .A2(_04251_),
    .B1(_04319_),
    .C1(_04288_),
    .X(_04384_));
 sky130_fd_sc_hd__nand3_2 _11982_ (.A(_04382_),
    .B(_04383_),
    .C(_04384_),
    .Y(_04385_));
 sky130_fd_sc_hd__a21o_1 _11983_ (.A1(_04354_),
    .A2(_04355_),
    .B1(_04353_),
    .X(_04386_));
 sky130_fd_sc_hd__a21o_1 _11984_ (.A1(_04383_),
    .A2(_04384_),
    .B1(_04382_),
    .X(_04387_));
 sky130_fd_sc_hd__nand4_1 _11985_ (.A(_04357_),
    .B(_04385_),
    .C(_04386_),
    .D(_04387_),
    .Y(_04388_));
 sky130_fd_sc_hd__a22o_1 _11986_ (.A1(_04357_),
    .A2(_04386_),
    .B1(_04387_),
    .B2(_04385_),
    .X(_04390_));
 sky130_fd_sc_hd__and2b_1 _11987_ (.A_N(_04287_),
    .B(_04321_),
    .X(_04391_));
 sky130_fd_sc_hd__a21oi_1 _11988_ (.A1(_04388_),
    .A2(_04390_),
    .B1(_04391_),
    .Y(_04392_));
 sky130_fd_sc_hd__inv_2 _11989_ (.A(_03987_),
    .Y(_04393_));
 sky130_fd_sc_hd__o211ai_1 _11990_ (.A1(_04393_),
    .A2(_03988_),
    .B1(_00530_),
    .C1(_01958_),
    .Y(_04394_));
 sky130_fd_sc_hd__a211o_1 _11991_ (.A1(_00530_),
    .A2(_01958_),
    .B1(_04393_),
    .C1(_03988_),
    .X(_04395_));
 sky130_fd_sc_hd__nand2_2 _11992_ (.A(_04394_),
    .B(_04395_),
    .Y(_04396_));
 sky130_fd_sc_hd__and3_1 _11993_ (.A(_04388_),
    .B(_04391_),
    .C(_04390_),
    .X(_04397_));
 sky130_fd_sc_hd__or3_4 _11994_ (.A(_04392_),
    .B(_04396_),
    .C(_04397_),
    .X(_04398_));
 sky130_fd_sc_hd__o21ai_1 _11995_ (.A1(_04392_),
    .A2(_04397_),
    .B1(_04396_),
    .Y(_04399_));
 sky130_fd_sc_hd__and3_1 _11996_ (.A(_04328_),
    .B(_04398_),
    .C(_04399_),
    .X(_04401_));
 sky130_fd_sc_hd__a21oi_4 _11997_ (.A1(_04398_),
    .A2(_04399_),
    .B1(_04328_),
    .Y(_04402_));
 sky130_fd_sc_hd__nor2_4 _11998_ (.A(_04401_),
    .B(_04402_),
    .Y(_04403_));
 sky130_fd_sc_hd__nor2_2 _11999_ (.A(_03990_),
    .B(_03992_),
    .Y(_04404_));
 sky130_fd_sc_hd__and2_1 _12000_ (.A(_03990_),
    .B(_03992_),
    .X(_04405_));
 sky130_fd_sc_hd__nor2_1 _12001_ (.A(_04404_),
    .B(_04405_),
    .Y(_04406_));
 sky130_fd_sc_hd__and4_1 _12002_ (.A(_04357_),
    .B(_04385_),
    .C(_04386_),
    .D(_04387_),
    .X(_04407_));
 sky130_fd_sc_hd__and2b_1 _12003_ (.A_N(_04340_),
    .B(_04342_),
    .X(_04408_));
 sky130_fd_sc_hd__and4_1 _12004_ (.A(_00257_),
    .B(_00670_),
    .C(_02090_),
    .D(_01780_),
    .X(_04409_));
 sky130_fd_sc_hd__a22oi_1 _12005_ (.A1(_00843_),
    .A2(_02090_),
    .B1(_02088_),
    .B2(_00844_),
    .Y(_04410_));
 sky130_fd_sc_hd__nor2_1 _12006_ (.A(_04409_),
    .B(_04410_),
    .Y(_04412_));
 sky130_fd_sc_hd__o21a_1 _12007_ (.A1(_04329_),
    .A2(_04333_),
    .B1(_04412_),
    .X(_04413_));
 sky130_fd_sc_hd__nor3_1 _12008_ (.A(_04329_),
    .B(_04333_),
    .C(_04412_),
    .Y(_04414_));
 sky130_fd_sc_hd__nor2_1 _12009_ (.A(_04413_),
    .B(_04414_),
    .Y(_04415_));
 sky130_fd_sc_hd__and2_1 _12010_ (.A(_04337_),
    .B(_04415_),
    .X(_04416_));
 sky130_fd_sc_hd__nor2_1 _12011_ (.A(_04337_),
    .B(_04415_),
    .Y(_04417_));
 sky130_fd_sc_hd__nor2_1 _12012_ (.A(_04416_),
    .B(_04417_),
    .Y(_04418_));
 sky130_fd_sc_hd__and2b_1 _12013_ (.A_N(_04408_),
    .B(_04418_),
    .X(_04419_));
 sky130_fd_sc_hd__and2b_1 _12014_ (.A_N(_04418_),
    .B(_04408_),
    .X(_04420_));
 sky130_fd_sc_hd__nor2_1 _12015_ (.A(_04419_),
    .B(_04420_),
    .Y(_04421_));
 sky130_fd_sc_hd__or2_1 _12016_ (.A(_04421_),
    .B(_04346_),
    .X(_04423_));
 sky130_fd_sc_hd__nand2_1 _12017_ (.A(_04421_),
    .B(_04346_),
    .Y(_04424_));
 sky130_fd_sc_hd__nand2_1 _12018_ (.A(_04423_),
    .B(_04424_),
    .Y(_04425_));
 sky130_fd_sc_hd__a31o_1 _12019_ (.A1(_04353_),
    .A2(_04354_),
    .A3(_04355_),
    .B1(_04351_),
    .X(_04426_));
 sky130_fd_sc_hd__xnor2_2 _12020_ (.A(_04425_),
    .B(_04426_),
    .Y(_04427_));
 sky130_fd_sc_hd__and2b_1 _12021_ (.A_N(_04369_),
    .B(_04371_),
    .X(_04428_));
 sky130_fd_sc_hd__and4_1 _12022_ (.A(_06626_),
    .B(_06450_),
    .C(_03683_),
    .D(_03679_),
    .X(_04429_));
 sky130_fd_sc_hd__a22oi_1 _12023_ (.A1(_06626_),
    .A2(_03683_),
    .B1(_03679_),
    .B2(_06450_),
    .Y(_04430_));
 sky130_fd_sc_hd__nor2_1 _12024_ (.A(_04429_),
    .B(_04430_),
    .Y(_04431_));
 sky130_fd_sc_hd__o21a_1 _12025_ (.A1(_04358_),
    .A2(_04362_),
    .B1(_04431_),
    .X(_04432_));
 sky130_fd_sc_hd__nor3_1 _12026_ (.A(_04358_),
    .B(_04362_),
    .C(_04431_),
    .Y(_04434_));
 sky130_fd_sc_hd__nor2_1 _12027_ (.A(_04432_),
    .B(_04434_),
    .Y(_04435_));
 sky130_fd_sc_hd__and2_1 _12028_ (.A(_04365_),
    .B(_04435_),
    .X(_04436_));
 sky130_fd_sc_hd__nor2_1 _12029_ (.A(_04365_),
    .B(_04435_),
    .Y(_04437_));
 sky130_fd_sc_hd__nor2_1 _12030_ (.A(_04436_),
    .B(_04437_),
    .Y(_04438_));
 sky130_fd_sc_hd__and2b_1 _12031_ (.A_N(_04428_),
    .B(_04438_),
    .X(_04439_));
 sky130_fd_sc_hd__and2b_1 _12032_ (.A_N(_04438_),
    .B(_04428_),
    .X(_04440_));
 sky130_fd_sc_hd__nor2_1 _12033_ (.A(_04439_),
    .B(_04440_),
    .Y(_04441_));
 sky130_fd_sc_hd__or2_1 _12034_ (.A(_04441_),
    .B(_04374_),
    .X(_04442_));
 sky130_fd_sc_hd__nand2_1 _12035_ (.A(_04441_),
    .B(_04374_),
    .Y(_04443_));
 sky130_fd_sc_hd__nand2_1 _12036_ (.A(_04442_),
    .B(_04443_),
    .Y(_04445_));
 sky130_fd_sc_hd__a31o_1 _12037_ (.A1(_04382_),
    .A2(_04383_),
    .A3(_04384_),
    .B1(_04380_),
    .X(_04446_));
 sky130_fd_sc_hd__xnor2_2 _12038_ (.A(_04445_),
    .B(_04446_),
    .Y(_04447_));
 sky130_fd_sc_hd__xor2_2 _12039_ (.A(_04427_),
    .B(_04447_),
    .X(_04448_));
 sky130_fd_sc_hd__xnor2_1 _12040_ (.A(_04407_),
    .B(_04448_),
    .Y(_04449_));
 sky130_fd_sc_hd__a21o_1 _12041_ (.A1(_04407_),
    .A2(_04448_),
    .B1(_04406_),
    .X(_04450_));
 sky130_fd_sc_hd__nor2_1 _12042_ (.A(_04407_),
    .B(_04448_),
    .Y(_04451_));
 sky130_fd_sc_hd__o2bb2a_2 _12043_ (.A1_N(_04406_),
    .A2_N(_04449_),
    .B1(_04450_),
    .B2(_04451_),
    .X(_04452_));
 sky130_fd_sc_hd__o21bai_4 _12044_ (.A1(_04396_),
    .A2(_04397_),
    .B1_N(_04392_),
    .Y(_04453_));
 sky130_fd_sc_hd__xor2_4 _12045_ (.A(_04452_),
    .B(_04453_),
    .X(_04454_));
 sky130_fd_sc_hd__xor2_1 _12046_ (.A(_04253_),
    .B(_04322_),
    .X(_04456_));
 sky130_fd_sc_hd__xnor2_1 _12047_ (.A(_04326_),
    .B(_04456_),
    .Y(_04457_));
 sky130_fd_sc_hd__xnor2_2 _12048_ (.A(_04142_),
    .B(_04252_),
    .Y(_04458_));
 sky130_fd_sc_hd__and3_1 _12049_ (.A(_04134_),
    .B(_04137_),
    .C(_04139_),
    .X(_04459_));
 sky130_fd_sc_hd__a21oi_1 _12050_ (.A1(_04137_),
    .A2(_04139_),
    .B1(_04134_),
    .Y(_04460_));
 sky130_fd_sc_hd__nor2_1 _12051_ (.A(_04459_),
    .B(_04460_),
    .Y(_04461_));
 sky130_fd_sc_hd__and3_1 _12052_ (.A(_04244_),
    .B(_04247_),
    .C(_04249_),
    .X(_04462_));
 sky130_fd_sc_hd__a21oi_1 _12053_ (.A1(_04247_),
    .A2(_04249_),
    .B1(_04244_),
    .Y(_04463_));
 sky130_fd_sc_hd__nor2_1 _12054_ (.A(_04462_),
    .B(_04463_),
    .Y(_04464_));
 sky130_fd_sc_hd__nand2_2 _12055_ (.A(_04461_),
    .B(_04464_),
    .Y(_04465_));
 sky130_fd_sc_hd__xnor2_1 _12056_ (.A(_03928_),
    .B(_03929_),
    .Y(_04467_));
 sky130_fd_sc_hd__a21boi_1 _12057_ (.A1(_04458_),
    .A2(_04465_),
    .B1_N(_04467_),
    .Y(_04468_));
 sky130_fd_sc_hd__o21ba_1 _12058_ (.A1(_04458_),
    .A2(_04465_),
    .B1_N(_04468_),
    .X(_04469_));
 sky130_fd_sc_hd__inv_2 _12059_ (.A(_04469_),
    .Y(_04470_));
 sky130_fd_sc_hd__and2_1 _12060_ (.A(_04457_),
    .B(_04470_),
    .X(_04471_));
 sky130_fd_sc_hd__xor2_1 _12061_ (.A(_04458_),
    .B(_04465_),
    .X(_04472_));
 sky130_fd_sc_hd__xnor2_1 _12062_ (.A(_04467_),
    .B(_04472_),
    .Y(_04473_));
 sky130_fd_sc_hd__or2_1 _12063_ (.A(_04461_),
    .B(_04464_),
    .X(_04474_));
 sky130_fd_sc_hd__xor2_1 _12064_ (.A(_04137_),
    .B(_04139_),
    .X(_04475_));
 sky130_fd_sc_hd__xor2_1 _12065_ (.A(_04247_),
    .B(_04249_),
    .X(_04476_));
 sky130_fd_sc_hd__and2_1 _12066_ (.A(_04475_),
    .B(_04476_),
    .X(_04478_));
 sky130_fd_sc_hd__a21o_1 _12067_ (.A1(_04465_),
    .A2(_04474_),
    .B1(_04478_),
    .X(_04479_));
 sky130_fd_sc_hd__a22oi_1 _12068_ (.A1(_03554_),
    .A2(_01183_),
    .B1(_01252_),
    .B2(_00530_),
    .Y(_04480_));
 sky130_fd_sc_hd__nor2_1 _12069_ (.A(_03929_),
    .B(_04480_),
    .Y(_04481_));
 sky130_fd_sc_hd__and3_1 _12070_ (.A(_04465_),
    .B(_04474_),
    .C(_04478_),
    .X(_04482_));
 sky130_fd_sc_hd__a21oi_1 _12071_ (.A1(_04479_),
    .A2(_04481_),
    .B1(_04482_),
    .Y(_04483_));
 sky130_fd_sc_hd__nor2_1 _12072_ (.A(_04473_),
    .B(_04483_),
    .Y(_04484_));
 sky130_fd_sc_hd__nor2_1 _12073_ (.A(_04457_),
    .B(_04470_),
    .Y(_04485_));
 sky130_fd_sc_hd__o21ba_1 _12074_ (.A1(_04471_),
    .A2(_04484_),
    .B1_N(_04485_),
    .X(_04486_));
 sky130_fd_sc_hd__nor2_1 _12075_ (.A(_04452_),
    .B(_04453_),
    .Y(_04487_));
 sky130_fd_sc_hd__nand2_1 _12076_ (.A(_04452_),
    .B(_04453_),
    .Y(_04489_));
 sky130_fd_sc_hd__o21a_1 _12077_ (.A1(_04487_),
    .A2(_04402_),
    .B1(_04489_),
    .X(_04490_));
 sky130_fd_sc_hd__a31oi_2 _12078_ (.A1(_04403_),
    .A2(_04454_),
    .A3(_04486_),
    .B1(_04490_),
    .Y(_04491_));
 sky130_fd_sc_hd__xnor2_4 _12079_ (.A(_03984_),
    .B(_04404_),
    .Y(_04492_));
 sky130_fd_sc_hd__and3_1 _12080_ (.A(_02246_),
    .B(_02426_),
    .C(_04330_),
    .X(_04493_));
 sky130_fd_sc_hd__and2_1 _12081_ (.A(_04413_),
    .B(_04493_),
    .X(_04494_));
 sky130_fd_sc_hd__nor2_1 _12082_ (.A(_04413_),
    .B(_04493_),
    .Y(_04495_));
 sky130_fd_sc_hd__nor2_1 _12083_ (.A(_04494_),
    .B(_04495_),
    .Y(_04496_));
 sky130_fd_sc_hd__o21a_1 _12084_ (.A1(_04416_),
    .A2(_04419_),
    .B1(_04496_),
    .X(_04497_));
 sky130_fd_sc_hd__nor3_1 _12085_ (.A(_04496_),
    .B(_04416_),
    .C(_04419_),
    .Y(_04498_));
 sky130_fd_sc_hd__nor2_2 _12086_ (.A(_04497_),
    .B(_04498_),
    .Y(_04500_));
 sky130_fd_sc_hd__o21a_1 _12087_ (.A1(_04346_),
    .A2(_04351_),
    .B1(_04421_),
    .X(_04501_));
 sky130_fd_sc_hd__a41o_2 _12088_ (.A1(_04353_),
    .A2(_04354_),
    .A3(_04355_),
    .A4(_04423_),
    .B1(_04501_),
    .X(_04502_));
 sky130_fd_sc_hd__xor2_2 _12089_ (.A(_04500_),
    .B(_04502_),
    .X(_04503_));
 sky130_fd_sc_hd__and3_1 _12090_ (.A(_06626_),
    .B(_03680_),
    .C(_04359_),
    .X(_04504_));
 sky130_fd_sc_hd__and2_1 _12091_ (.A(_04432_),
    .B(_04504_),
    .X(_04505_));
 sky130_fd_sc_hd__nor2_1 _12092_ (.A(_04432_),
    .B(_04504_),
    .Y(_04506_));
 sky130_fd_sc_hd__nor2_1 _12093_ (.A(_04505_),
    .B(_04506_),
    .Y(_04507_));
 sky130_fd_sc_hd__o21a_1 _12094_ (.A1(_04436_),
    .A2(_04439_),
    .B1(_04507_),
    .X(_04508_));
 sky130_fd_sc_hd__nor3_1 _12095_ (.A(_04507_),
    .B(_04436_),
    .C(_04439_),
    .Y(_04509_));
 sky130_fd_sc_hd__nor2_2 _12096_ (.A(_04508_),
    .B(_04509_),
    .Y(_04511_));
 sky130_fd_sc_hd__o21a_1 _12097_ (.A1(_04374_),
    .A2(_04380_),
    .B1(_04441_),
    .X(_04512_));
 sky130_fd_sc_hd__a41o_2 _12098_ (.A1(_04382_),
    .A2(_04383_),
    .A3(_04384_),
    .A4(_04442_),
    .B1(_04512_),
    .X(_04513_));
 sky130_fd_sc_hd__xor2_2 _12099_ (.A(_04511_),
    .B(_04513_),
    .X(_04514_));
 sky130_fd_sc_hd__xnor2_2 _12100_ (.A(_04503_),
    .B(_04514_),
    .Y(_04515_));
 sky130_fd_sc_hd__nand2_1 _12101_ (.A(_04427_),
    .B(_04447_),
    .Y(_04516_));
 sky130_fd_sc_hd__nand2_1 _12102_ (.A(_04515_),
    .B(_04516_),
    .Y(_04517_));
 sky130_fd_sc_hd__nor2_1 _12103_ (.A(_04515_),
    .B(_04516_),
    .Y(_04518_));
 sky130_fd_sc_hd__a21o_2 _12104_ (.A1(_04492_),
    .A2(_04517_),
    .B1(_04518_),
    .X(_04519_));
 sky130_fd_sc_hd__and3_1 _12105_ (.A(_03996_),
    .B(_03983_),
    .C(_03994_),
    .X(_04520_));
 sky130_fd_sc_hd__nor2_2 _12106_ (.A(_03997_),
    .B(_04520_),
    .Y(_04522_));
 sky130_fd_sc_hd__and2_2 _12107_ (.A(_04503_),
    .B(_04514_),
    .X(_04523_));
 sky130_fd_sc_hd__or3_1 _12108_ (.A(_04409_),
    .B(_04494_),
    .C(_04497_),
    .X(_04524_));
 sky130_fd_sc_hd__a21oi_4 _12109_ (.A1(_04500_),
    .A2(_04502_),
    .B1(_04524_),
    .Y(_04525_));
 sky130_fd_sc_hd__or3_1 _12110_ (.A(_04429_),
    .B(_04505_),
    .C(_04508_),
    .X(_04526_));
 sky130_fd_sc_hd__a21oi_4 _12111_ (.A1(_04511_),
    .A2(_04513_),
    .B1(_04526_),
    .Y(_04527_));
 sky130_fd_sc_hd__xor2_4 _12112_ (.A(_04525_),
    .B(_04527_),
    .X(_04528_));
 sky130_fd_sc_hd__xnor2_2 _12113_ (.A(_04523_),
    .B(_04528_),
    .Y(_04529_));
 sky130_fd_sc_hd__xnor2_4 _12114_ (.A(_04522_),
    .B(_04529_),
    .Y(_04530_));
 sky130_fd_sc_hd__xor2_4 _12115_ (.A(_04519_),
    .B(_04530_),
    .X(_04531_));
 sky130_fd_sc_hd__xnor2_2 _12116_ (.A(_04515_),
    .B(_04516_),
    .Y(_04533_));
 sky130_fd_sc_hd__xnor2_4 _12117_ (.A(_04492_),
    .B(_04533_),
    .Y(_04534_));
 sky130_fd_sc_hd__and2b_2 _12118_ (.A_N(_04451_),
    .B(_04450_),
    .X(_04535_));
 sky130_fd_sc_hd__xor2_4 _12119_ (.A(_04534_),
    .B(_04535_),
    .X(_04536_));
 sky130_fd_sc_hd__nand2_1 _12120_ (.A(_04531_),
    .B(_04536_),
    .Y(_04537_));
 sky130_fd_sc_hd__and2_1 _12121_ (.A(_03956_),
    .B(_04001_),
    .X(_04538_));
 sky130_fd_sc_hd__nor2_1 _12122_ (.A(_04002_),
    .B(_04538_),
    .Y(_04539_));
 sky130_fd_sc_hd__inv_2 _12123_ (.A(_04539_),
    .Y(_04540_));
 sky130_fd_sc_hd__nor2_1 _12124_ (.A(_04525_),
    .B(_04527_),
    .Y(_04541_));
 sky130_fd_sc_hd__or3_1 _12125_ (.A(_04000_),
    .B(_03969_),
    .C(_03997_),
    .X(_04542_));
 sky130_fd_sc_hd__and2_1 _12126_ (.A(_04001_),
    .B(_04542_),
    .X(_04544_));
 sky130_fd_sc_hd__and2_1 _12127_ (.A(_04541_),
    .B(_04544_),
    .X(_04545_));
 sky130_fd_sc_hd__mux2_2 _12128_ (.A0(_04540_),
    .A1(_03955_),
    .S(_04545_),
    .X(_04546_));
 sky130_fd_sc_hd__nor2_1 _12129_ (.A(_04541_),
    .B(_04544_),
    .Y(_04547_));
 sky130_fd_sc_hd__or2_4 _12130_ (.A(_04545_),
    .B(_04547_),
    .X(_04548_));
 sky130_fd_sc_hd__a21o_1 _12131_ (.A1(_04523_),
    .A2(_04528_),
    .B1(_04522_),
    .X(_04549_));
 sky130_fd_sc_hd__o21ai_4 _12132_ (.A1(_04523_),
    .A2(_04528_),
    .B1(_04549_),
    .Y(_04550_));
 sky130_fd_sc_hd__xor2_4 _12133_ (.A(_04548_),
    .B(_04550_),
    .X(_04551_));
 sky130_fd_sc_hd__or2b_1 _12134_ (.A(_04546_),
    .B_N(_04551_),
    .X(_04552_));
 sky130_fd_sc_hd__nor2_1 _12135_ (.A(_04537_),
    .B(_04552_),
    .Y(_04553_));
 sky130_fd_sc_hd__and2b_1 _12136_ (.A_N(_04491_),
    .B(_04553_),
    .X(_04555_));
 sky130_fd_sc_hd__and2b_1 _12137_ (.A_N(_04482_),
    .B(_04479_),
    .X(_04556_));
 sky130_fd_sc_hd__xnor2_1 _12138_ (.A(_04481_),
    .B(_04556_),
    .Y(_04557_));
 sky130_fd_sc_hd__nor2_1 _12139_ (.A(_02596_),
    .B(_02644_),
    .Y(_04558_));
 sky130_fd_sc_hd__a21oi_2 _12140_ (.A1(_02596_),
    .A2(_02644_),
    .B1(_02693_),
    .Y(_04559_));
 sky130_fd_sc_hd__nor2_1 _12141_ (.A(_04475_),
    .B(_04476_),
    .Y(_04560_));
 sky130_fd_sc_hd__or2_1 _12142_ (.A(_04478_),
    .B(_04560_),
    .X(_04561_));
 sky130_fd_sc_hd__o21a_1 _12143_ (.A1(_04558_),
    .A2(_04559_),
    .B1(_04561_),
    .X(_04562_));
 sky130_fd_sc_hd__nand2_1 _12144_ (.A(_00530_),
    .B(_01183_),
    .Y(_04563_));
 sky130_fd_sc_hd__o31a_1 _12145_ (.A1(_04558_),
    .A2(_04561_),
    .A3(_04559_),
    .B1(_04563_),
    .X(_04564_));
 sky130_fd_sc_hd__nor3_2 _12146_ (.A(_04557_),
    .B(_04562_),
    .C(_04564_),
    .Y(_04566_));
 sky130_fd_sc_hd__inv_2 _12147_ (.A(_04566_),
    .Y(_04567_));
 sky130_fd_sc_hd__o21ai_1 _12148_ (.A1(_04558_),
    .A2(_04559_),
    .B1(_04561_),
    .Y(_04568_));
 sky130_fd_sc_hd__or3_1 _12149_ (.A(_04558_),
    .B(_04561_),
    .C(_04559_),
    .X(_04569_));
 sky130_fd_sc_hd__a21o_1 _12150_ (.A1(_04568_),
    .A2(_04569_),
    .B1(_04563_),
    .X(_04570_));
 sky130_fd_sc_hd__nand3_2 _12151_ (.A(_04568_),
    .B(_04563_),
    .C(_04569_),
    .Y(_04571_));
 sky130_fd_sc_hd__nand2_1 _12152_ (.A(_02694_),
    .B(_02698_),
    .Y(_04572_));
 sky130_fd_sc_hd__a21o_1 _12153_ (.A1(_04570_),
    .A2(_04571_),
    .B1(_04572_),
    .X(_04573_));
 sky130_fd_sc_hd__o21a_1 _12154_ (.A1(_04562_),
    .A2(_04564_),
    .B1(_04557_),
    .X(_04574_));
 sky130_fd_sc_hd__a21oi_4 _12155_ (.A1(_04567_),
    .A2(_04573_),
    .B1(_04574_),
    .Y(_04575_));
 sky130_fd_sc_hd__inv_2 _12156_ (.A(_02699_),
    .Y(_04577_));
 sky130_fd_sc_hd__nor2_2 _12157_ (.A(_04566_),
    .B(_04574_),
    .Y(_04578_));
 sky130_fd_sc_hd__nand2_1 _12158_ (.A(_04570_),
    .B(_04571_),
    .Y(_04579_));
 sky130_fd_sc_hd__o2111a_4 _12159_ (.A1(_02476_),
    .A2(_02480_),
    .B1(_04577_),
    .C1(_04578_),
    .D1(_04579_),
    .X(_04580_));
 sky130_fd_sc_hd__nor2_4 _12160_ (.A(_04471_),
    .B(_04485_),
    .Y(_04581_));
 sky130_fd_sc_hd__nand2_1 _12161_ (.A(_04473_),
    .B(_04483_),
    .Y(_04582_));
 sky130_fd_sc_hd__or2b_1 _12162_ (.A(_04484_),
    .B_N(_04582_),
    .X(_04583_));
 sky130_fd_sc_hd__inv_2 _12163_ (.A(_04583_),
    .Y(_04584_));
 sky130_fd_sc_hd__and4_1 _12164_ (.A(_04581_),
    .B(_04584_),
    .C(_04403_),
    .D(_04454_),
    .X(_04585_));
 sky130_fd_sc_hd__o211a_1 _12165_ (.A1(_04575_),
    .A2(_04580_),
    .B1(_04585_),
    .C1(_04553_),
    .X(_04586_));
 sky130_fd_sc_hd__and2_1 _12166_ (.A(_04519_),
    .B(_04530_),
    .X(_04588_));
 sky130_fd_sc_hd__and2_1 _12167_ (.A(_04534_),
    .B(_04535_),
    .X(_04589_));
 sky130_fd_sc_hd__nor2_1 _12168_ (.A(_04519_),
    .B(_04530_),
    .Y(_04590_));
 sky130_fd_sc_hd__o21bai_1 _12169_ (.A1(_04588_),
    .A2(_04589_),
    .B1_N(_04590_),
    .Y(_04591_));
 sky130_fd_sc_hd__nor2_1 _12170_ (.A(_04548_),
    .B(_04550_),
    .Y(_04592_));
 sky130_fd_sc_hd__o21ai_1 _12171_ (.A1(_04545_),
    .A2(_04592_),
    .B1(_04539_),
    .Y(_04593_));
 sky130_fd_sc_hd__o21ai_1 _12172_ (.A1(_04591_),
    .A2(_04552_),
    .B1(_04593_),
    .Y(_04594_));
 sky130_fd_sc_hd__or3_4 _12173_ (.A(_04555_),
    .B(_04586_),
    .C(_04594_),
    .X(_04595_));
 sky130_fd_sc_hd__or4b_4 _12174_ (.A(_04025_),
    .B(_04028_),
    .C(_04032_),
    .D_N(_04595_),
    .X(_04596_));
 sky130_fd_sc_hd__a211oi_1 _12175_ (.A1(_03728_),
    .A2(_04017_),
    .B1(_04021_),
    .C1(_03725_),
    .Y(_04597_));
 sky130_fd_sc_hd__nand2_1 _12176_ (.A(_04018_),
    .B(_04019_),
    .Y(_04599_));
 sky130_fd_sc_hd__o211a_4 _12177_ (.A1(_04024_),
    .A2(net186),
    .B1(_04597_),
    .C1(_04599_),
    .X(_04600_));
 sky130_fd_sc_hd__xor2_2 _12178_ (.A(_03677_),
    .B(_04600_),
    .X(_04601_));
 sky130_fd_sc_hd__a21o_1 _12179_ (.A1(_03589_),
    .A2(_03551_),
    .B1(_03583_),
    .X(_04602_));
 sky130_fd_sc_hd__or2_2 _12180_ (.A(_03582_),
    .B(_03583_),
    .X(_04603_));
 sky130_fd_sc_hd__and2_1 _12181_ (.A(_03548_),
    .B(_03549_),
    .X(_04604_));
 sky130_fd_sc_hd__xnor2_1 _12182_ (.A(_03550_),
    .B(_04604_),
    .Y(_04605_));
 sky130_fd_sc_hd__a2111o_2 _12183_ (.A1(_02382_),
    .A2(_02385_),
    .B1(_02588_),
    .C1(_04603_),
    .D1(_04605_),
    .X(_04606_));
 sky130_fd_sc_hd__or3b_1 _12184_ (.A(_03608_),
    .B(_03578_),
    .C_N(_03610_),
    .X(_04607_));
 sky130_fd_sc_hd__nand2_1 _12185_ (.A(_03614_),
    .B(_03602_),
    .Y(_04608_));
 sky130_fd_sc_hd__a211o_1 _12186_ (.A1(_04602_),
    .A2(_04606_),
    .B1(_04607_),
    .C1(_04608_),
    .X(_04610_));
 sky130_fd_sc_hd__nand2_1 _12187_ (.A(_03613_),
    .B(_03623_),
    .Y(_04611_));
 sky130_fd_sc_hd__or2b_1 _12188_ (.A(_03493_),
    .B_N(_03622_),
    .X(_04612_));
 sky130_fd_sc_hd__or2_1 _12189_ (.A(_04611_),
    .B(_04612_),
    .X(_04613_));
 sky130_fd_sc_hd__o21ai_1 _12190_ (.A1(_03608_),
    .A2(_03575_),
    .B1(_03610_),
    .Y(_04614_));
 sky130_fd_sc_hd__or2b_1 _12191_ (.A(_03533_),
    .B_N(_03514_),
    .X(_04615_));
 sky130_fd_sc_hd__o21a_1 _12192_ (.A1(_03534_),
    .A2(_03617_),
    .B1(_04615_),
    .X(_04616_));
 sky130_fd_sc_hd__o21ba_1 _12193_ (.A1(_04614_),
    .A2(_04608_),
    .B1_N(_04616_),
    .X(_04617_));
 sky130_fd_sc_hd__or2_1 _12194_ (.A(_04617_),
    .B(_04613_),
    .X(_04618_));
 sky130_fd_sc_hd__or2_1 _12195_ (.A(_03484_),
    .B(_03486_),
    .X(_04619_));
 sky130_fd_sc_hd__o21ai_1 _12196_ (.A1(_03487_),
    .A2(_03512_),
    .B1(_04619_),
    .Y(_04621_));
 sky130_fd_sc_hd__o21ai_1 _12197_ (.A1(_03453_),
    .A2(_03468_),
    .B1(_03492_),
    .Y(_04622_));
 sky130_fd_sc_hd__o21a_1 _12198_ (.A1(_04621_),
    .A2(_04612_),
    .B1(_04622_),
    .X(_04623_));
 sky130_fd_sc_hd__o211ai_4 _12199_ (.A1(_04610_),
    .A2(_04613_),
    .B1(_04618_),
    .C1(_04623_),
    .Y(_04624_));
 sky130_fd_sc_hd__or3b_1 _12200_ (.A(_03053_),
    .B(_03673_),
    .C_N(_04624_),
    .X(_04625_));
 sky130_fd_sc_hd__xor2_2 _12201_ (.A(_03667_),
    .B(_04625_),
    .X(_04626_));
 sky130_fd_sc_hd__xnor2_4 _12202_ (.A(_04024_),
    .B(_04596_),
    .Y(_04627_));
 sky130_fd_sc_hd__or2_1 _12203_ (.A(_04626_),
    .B(_04627_),
    .X(_04628_));
 sky130_fd_sc_hd__nor2_1 _12204_ (.A(_04601_),
    .B(_04628_),
    .Y(_04629_));
 sky130_fd_sc_hd__and4_1 _12205_ (.A(_00374_),
    .B(_00784_),
    .C(_01953_),
    .D(_02134_),
    .X(_04630_));
 sky130_fd_sc_hd__a22o_1 _12206_ (.A1(_00784_),
    .A2(_01953_),
    .B1(_02134_),
    .B2(_00374_),
    .X(_04632_));
 sky130_fd_sc_hd__and4b_1 _12207_ (.A_N(_04630_),
    .B(_03682_),
    .C(_00379_),
    .D(_04632_),
    .X(_04633_));
 sky130_fd_sc_hd__a22oi_1 _12208_ (.A1(_01518_),
    .A2(_01954_),
    .B1(_02135_),
    .B2(_00375_),
    .Y(_04634_));
 sky130_fd_sc_hd__o2bb2a_1 _12209_ (.A1_N(_00379_),
    .A2_N(_03682_),
    .B1(_04634_),
    .B2(_04630_),
    .X(_04635_));
 sky130_fd_sc_hd__or2_1 _12210_ (.A(_04633_),
    .B(_04635_),
    .X(_04636_));
 sky130_fd_sc_hd__and4_1 _12211_ (.A(_00376_),
    .B(_00379_),
    .C(_01954_),
    .D(_02135_),
    .X(_04637_));
 sky130_fd_sc_hd__xnor2_1 _12212_ (.A(_04636_),
    .B(_04637_),
    .Y(_04638_));
 sky130_fd_sc_hd__and4_1 _12213_ (.A(_00605_),
    .B(_01507_),
    .C(_01179_),
    .D(_01254_),
    .X(_04639_));
 sky130_fd_sc_hd__a22o_1 _12214_ (.A1(_01507_),
    .A2(_01179_),
    .B1(_01254_),
    .B2(_00605_),
    .X(_04640_));
 sky130_fd_sc_hd__and4b_1 _12215_ (.A_N(_04639_),
    .B(_03750_),
    .C(_00458_),
    .D(_04640_),
    .X(_04641_));
 sky130_fd_sc_hd__a22oi_1 _12216_ (.A1(_01664_),
    .A2(_01180_),
    .B1(_01249_),
    .B2(_00607_),
    .Y(_04643_));
 sky130_fd_sc_hd__o2bb2a_1 _12217_ (.A1_N(_00458_),
    .A2_N(_03750_),
    .B1(_04643_),
    .B2(_04639_),
    .X(_04644_));
 sky130_fd_sc_hd__or2_1 _12218_ (.A(_04641_),
    .B(_04644_),
    .X(_04645_));
 sky130_fd_sc_hd__nand4_4 _12219_ (.A(_00459_),
    .B(_00608_),
    .C(_01180_),
    .D(_01249_),
    .Y(_04646_));
 sky130_fd_sc_hd__nor2_1 _12220_ (.A(_04645_),
    .B(_04646_),
    .Y(_04647_));
 sky130_fd_sc_hd__and2_1 _12221_ (.A(_04645_),
    .B(_04646_),
    .X(_04648_));
 sky130_fd_sc_hd__or2_1 _12222_ (.A(_04647_),
    .B(_04648_),
    .X(_04649_));
 sky130_fd_sc_hd__a22o_1 _12223_ (.A1(_00778_),
    .A2(_01248_),
    .B1(_02117_),
    .B2(_00783_),
    .X(_04650_));
 sky130_fd_sc_hd__and4_1 _12224_ (.A(_00783_),
    .B(_00778_),
    .C(_01248_),
    .D(_02117_),
    .X(_04651_));
 sky130_fd_sc_hd__a31o_1 _12225_ (.A1(_00375_),
    .A2(_03744_),
    .A3(_04650_),
    .B1(_04651_),
    .X(_04652_));
 sky130_fd_sc_hd__nand4_2 _12226_ (.A(_01518_),
    .B(_01517_),
    .C(_03738_),
    .D(_03744_),
    .Y(_04654_));
 sky130_fd_sc_hd__a22o_1 _12227_ (.A1(_01517_),
    .A2(_03738_),
    .B1(_03744_),
    .B2(_01518_),
    .X(_04655_));
 sky130_fd_sc_hd__and3_1 _12228_ (.A(_04652_),
    .B(_04654_),
    .C(_04655_),
    .X(_04656_));
 sky130_fd_sc_hd__nand2_1 _12229_ (.A(_01518_),
    .B(_03750_),
    .Y(_04657_));
 sky130_fd_sc_hd__and3_1 _12230_ (.A(_01517_),
    .B(_03748_),
    .C(_04657_),
    .X(_04658_));
 sky130_fd_sc_hd__nand2_1 _12231_ (.A(_04656_),
    .B(_04658_),
    .Y(_04659_));
 sky130_fd_sc_hd__or2_1 _12232_ (.A(_04656_),
    .B(_04658_),
    .X(_04660_));
 sky130_fd_sc_hd__nand2_1 _12233_ (.A(_04659_),
    .B(_04660_),
    .Y(_04661_));
 sky130_fd_sc_hd__a22o_1 _12234_ (.A1(_00778_),
    .A2(_01178_),
    .B1(_01248_),
    .B2(_00783_),
    .X(_04662_));
 sky130_fd_sc_hd__and4_1 _12235_ (.A(_00783_),
    .B(_00778_),
    .C(_01178_),
    .D(_01248_),
    .X(_04663_));
 sky130_fd_sc_hd__a31o_1 _12236_ (.A1(_00375_),
    .A2(_03750_),
    .A3(_04662_),
    .B1(_04663_),
    .X(_04665_));
 sky130_fd_sc_hd__and2b_1 _12237_ (.A_N(_04651_),
    .B(_04650_),
    .X(_04666_));
 sky130_fd_sc_hd__nand2_1 _12238_ (.A(_00375_),
    .B(_02120_),
    .Y(_04667_));
 sky130_fd_sc_hd__xnor2_2 _12239_ (.A(_04666_),
    .B(_04667_),
    .Y(_04668_));
 sky130_fd_sc_hd__a21oi_1 _12240_ (.A1(_04654_),
    .A2(_04655_),
    .B1(_04652_),
    .Y(_04669_));
 sky130_fd_sc_hd__nor2_1 _12241_ (.A(_04656_),
    .B(_04669_),
    .Y(_04670_));
 sky130_fd_sc_hd__and3_1 _12242_ (.A(_04665_),
    .B(_04668_),
    .C(_04670_),
    .X(_04671_));
 sky130_fd_sc_hd__a21oi_1 _12243_ (.A1(_04665_),
    .A2(_04668_),
    .B1(_04670_),
    .Y(_04672_));
 sky130_fd_sc_hd__nor2_1 _12244_ (.A(_04671_),
    .B(_04672_),
    .Y(_04673_));
 sky130_fd_sc_hd__a22o_1 _12245_ (.A1(_00783_),
    .A2(_01178_),
    .B1(_01248_),
    .B2(_04037_),
    .X(_04674_));
 sky130_fd_sc_hd__and4_1 _12246_ (.A(_04037_),
    .B(_00783_),
    .C(_01178_),
    .D(_01248_),
    .X(_04676_));
 sky130_fd_sc_hd__a31o_1 _12247_ (.A1(_00378_),
    .A2(_02119_),
    .A3(_04674_),
    .B1(_04676_),
    .X(_04677_));
 sky130_fd_sc_hd__and3_1 _12248_ (.A(_00379_),
    .B(_03748_),
    .C(_04677_),
    .X(_04678_));
 sky130_fd_sc_hd__or2b_1 _12249_ (.A(_04663_),
    .B_N(_04662_),
    .X(_04679_));
 sky130_fd_sc_hd__nand2_1 _12250_ (.A(_00375_),
    .B(_03738_),
    .Y(_04680_));
 sky130_fd_sc_hd__xnor2_1 _12251_ (.A(_04679_),
    .B(_04680_),
    .Y(_04681_));
 sky130_fd_sc_hd__nand2_1 _12252_ (.A(_00378_),
    .B(_02120_),
    .Y(_04682_));
 sky130_fd_sc_hd__xnor2_1 _12253_ (.A(_04677_),
    .B(_04682_),
    .Y(_04683_));
 sky130_fd_sc_hd__and2b_1 _12254_ (.A_N(_04681_),
    .B(_04683_),
    .X(_04684_));
 sky130_fd_sc_hd__xor2_1 _12255_ (.A(_04665_),
    .B(_04668_),
    .X(_04685_));
 sky130_fd_sc_hd__or3_1 _12256_ (.A(_04678_),
    .B(_04684_),
    .C(_04685_),
    .X(_04687_));
 sky130_fd_sc_hd__or2b_2 _12257_ (.A(_04676_),
    .B_N(_04674_),
    .X(_04688_));
 sky130_fd_sc_hd__nand2_2 _12258_ (.A(_00378_),
    .B(_03738_),
    .Y(_04689_));
 sky130_fd_sc_hd__xnor2_4 _12259_ (.A(_04688_),
    .B(_04689_),
    .Y(_04690_));
 sky130_fd_sc_hd__and4_2 _12260_ (.A(_00376_),
    .B(_00378_),
    .C(_01180_),
    .D(_01249_),
    .X(_04691_));
 sky130_fd_sc_hd__and2b_1 _12261_ (.A_N(_04690_),
    .B(_04691_),
    .X(_04692_));
 sky130_fd_sc_hd__xnor2_1 _12262_ (.A(_04681_),
    .B(_04683_),
    .Y(_04693_));
 sky130_fd_sc_hd__and2_1 _12263_ (.A(_04692_),
    .B(_04693_),
    .X(_04694_));
 sky130_fd_sc_hd__o21a_1 _12264_ (.A1(_04678_),
    .A2(_04684_),
    .B1(_04685_),
    .X(_04695_));
 sky130_fd_sc_hd__a21o_1 _12265_ (.A1(_04687_),
    .A2(_04694_),
    .B1(_04695_),
    .X(_04696_));
 sky130_fd_sc_hd__a21o_1 _12266_ (.A1(_04673_),
    .A2(_04696_),
    .B1(_04671_),
    .X(_04698_));
 sky130_fd_sc_hd__xor2_2 _12267_ (.A(_04661_),
    .B(_04698_),
    .X(_04699_));
 sky130_fd_sc_hd__xor2_1 _12268_ (.A(_04649_),
    .B(_04699_),
    .X(_04700_));
 sky130_fd_sc_hd__xnor2_1 _12269_ (.A(_04638_),
    .B(_04700_),
    .Y(_04701_));
 sky130_fd_sc_hd__a22o_1 _12270_ (.A1(_03414_),
    .A2(_01181_),
    .B1(_01250_),
    .B2(_01066_),
    .X(_04702_));
 sky130_fd_sc_hd__a21oi_1 _12271_ (.A1(_04687_),
    .A2(_04694_),
    .B1(_04695_),
    .Y(_04703_));
 sky130_fd_sc_hd__xnor2_1 _12272_ (.A(_04673_),
    .B(_04703_),
    .Y(_04704_));
 sky130_fd_sc_hd__a21o_1 _12273_ (.A1(_04646_),
    .A2(_04702_),
    .B1(_04704_),
    .X(_04705_));
 sky130_fd_sc_hd__a22oi_1 _12274_ (.A1(_00376_),
    .A2(_01955_),
    .B1(_03686_),
    .B2(_00380_),
    .Y(_04706_));
 sky130_fd_sc_hd__nor2_1 _12275_ (.A(_04637_),
    .B(_04706_),
    .Y(_04707_));
 sky130_fd_sc_hd__nand3_1 _12276_ (.A(_04646_),
    .B(_04702_),
    .C(_04704_),
    .Y(_04709_));
 sky130_fd_sc_hd__a21bo_1 _12277_ (.A1(_04705_),
    .A2(_04707_),
    .B1_N(_04709_),
    .X(_04710_));
 sky130_fd_sc_hd__and2b_1 _12278_ (.A_N(_04701_),
    .B(_04710_),
    .X(_04711_));
 sky130_fd_sc_hd__or2b_1 _12279_ (.A(_04710_),
    .B_N(_04701_),
    .X(_04712_));
 sky130_fd_sc_hd__or2b_1 _12280_ (.A(_04711_),
    .B_N(_04712_),
    .X(_04713_));
 sky130_fd_sc_hd__clkbuf_4 _12281_ (.A(_01066_),
    .X(_04714_));
 sky130_fd_sc_hd__or2b_1 _12282_ (.A(_04695_),
    .B_N(_04687_),
    .X(_04715_));
 sky130_fd_sc_hd__xnor2_1 _12283_ (.A(_04715_),
    .B(_04694_),
    .Y(_04716_));
 sky130_fd_sc_hd__a21o_1 _12284_ (.A1(_04714_),
    .A2(_01182_),
    .B1(_04716_),
    .X(_04717_));
 sky130_fd_sc_hd__and3_1 _12285_ (.A(_04714_),
    .B(_01181_),
    .C(_04716_),
    .X(_04718_));
 sky130_fd_sc_hd__a21o_1 _12286_ (.A1(_00380_),
    .A2(_01956_),
    .B1(_04718_),
    .X(_04720_));
 sky130_fd_sc_hd__nand2_1 _12287_ (.A(_04717_),
    .B(_04720_),
    .Y(_04721_));
 sky130_fd_sc_hd__nand2_1 _12288_ (.A(_04709_),
    .B(_04705_),
    .Y(_04722_));
 sky130_fd_sc_hd__xor2_1 _12289_ (.A(_04707_),
    .B(_04722_),
    .X(_04723_));
 sky130_fd_sc_hd__nor2_1 _12290_ (.A(_04721_),
    .B(_04723_),
    .Y(_04724_));
 sky130_fd_sc_hd__xor2_2 _12291_ (.A(_04713_),
    .B(_04724_),
    .X(_04725_));
 sky130_fd_sc_hd__a22o_1 _12292_ (.A1(_02187_),
    .A2(_01601_),
    .B1(_02189_),
    .B2(_00575_),
    .X(_04726_));
 sky130_fd_sc_hd__and4_1 _12293_ (.A(_00575_),
    .B(_01664_),
    .C(_01601_),
    .D(_01505_),
    .X(_04727_));
 sky130_fd_sc_hd__a31o_1 _12294_ (.A1(_03414_),
    .A2(_02426_),
    .A3(_04726_),
    .B1(_04727_),
    .X(_04728_));
 sky130_fd_sc_hd__and4_1 _12295_ (.A(_02188_),
    .B(_02427_),
    .C(_02190_),
    .D(_02088_),
    .X(_04729_));
 sky130_fd_sc_hd__a22oi_1 _12296_ (.A1(_02427_),
    .A2(_02190_),
    .B1(_02088_),
    .B2(_02188_),
    .Y(_04731_));
 sky130_fd_sc_hd__nor2_1 _12297_ (.A(_04729_),
    .B(_04731_),
    .Y(_04732_));
 sky130_fd_sc_hd__and2_1 _12298_ (.A(_04728_),
    .B(_04732_),
    .X(_04733_));
 sky130_fd_sc_hd__nand2_1 _12299_ (.A(_02188_),
    .B(_02427_),
    .Y(_04734_));
 sky130_fd_sc_hd__and3_1 _12300_ (.A(_02190_),
    .B(_02426_),
    .C(_04734_),
    .X(_04735_));
 sky130_fd_sc_hd__xor2_2 _12301_ (.A(_04733_),
    .B(_04735_),
    .X(_04736_));
 sky130_fd_sc_hd__and4_1 _12302_ (.A(_00415_),
    .B(_00575_),
    .C(_01664_),
    .D(_01505_),
    .X(_04737_));
 sky130_fd_sc_hd__a22oi_1 _12303_ (.A1(_01288_),
    .A2(_02187_),
    .B1(_02189_),
    .B2(_00416_),
    .Y(_04738_));
 sky130_fd_sc_hd__and4bb_1 _12304_ (.A_N(_04737_),
    .B_N(_04738_),
    .C(_00608_),
    .D(_01601_),
    .X(_04739_));
 sky130_fd_sc_hd__and2b_1 _12305_ (.A_N(_04727_),
    .B(_04726_),
    .X(_04740_));
 sky130_fd_sc_hd__nand2_1 _12306_ (.A(_01400_),
    .B(_01780_),
    .Y(_04742_));
 sky130_fd_sc_hd__xnor2_1 _12307_ (.A(_04740_),
    .B(_04742_),
    .Y(_04743_));
 sky130_fd_sc_hd__o21a_1 _12308_ (.A1(_04737_),
    .A2(_04739_),
    .B1(_04743_),
    .X(_04744_));
 sky130_fd_sc_hd__nor2_1 _12309_ (.A(_04728_),
    .B(_04732_),
    .Y(_04745_));
 sky130_fd_sc_hd__nor2_1 _12310_ (.A(_04733_),
    .B(_04745_),
    .Y(_04746_));
 sky130_fd_sc_hd__a22o_1 _12311_ (.A1(_00607_),
    .A2(_00575_),
    .B1(_01664_),
    .B2(_00415_),
    .X(_04747_));
 sky130_fd_sc_hd__and3_1 _12312_ (.A(_00415_),
    .B(_00607_),
    .C(_01664_),
    .X(_04748_));
 sky130_fd_sc_hd__a32o_1 _12313_ (.A1(_00459_),
    .A2(_01601_),
    .A3(_04747_),
    .B1(_04748_),
    .B2(_01288_),
    .X(_04749_));
 sky130_fd_sc_hd__and3_1 _12314_ (.A(_00459_),
    .B(_01780_),
    .C(_04749_),
    .X(_04750_));
 sky130_fd_sc_hd__o2bb2a_1 _12315_ (.A1_N(_00608_),
    .A2_N(_01601_),
    .B1(_04737_),
    .B2(_04738_),
    .X(_04751_));
 sky130_fd_sc_hd__or2_1 _12316_ (.A(_04739_),
    .B(_04751_),
    .X(_04753_));
 sky130_fd_sc_hd__a21oi_1 _12317_ (.A1(_00460_),
    .A2(_02088_),
    .B1(_04749_),
    .Y(_04754_));
 sky130_fd_sc_hd__nor2_1 _12318_ (.A(_04750_),
    .B(_04754_),
    .Y(_04755_));
 sky130_fd_sc_hd__and2b_1 _12319_ (.A_N(_04753_),
    .B(_04755_),
    .X(_04756_));
 sky130_fd_sc_hd__nor3_1 _12320_ (.A(_04737_),
    .B(_04739_),
    .C(_04743_),
    .Y(_04757_));
 sky130_fd_sc_hd__nor2_1 _12321_ (.A(_04744_),
    .B(_04757_),
    .Y(_04758_));
 sky130_fd_sc_hd__o21ai_1 _12322_ (.A1(_04750_),
    .A2(_04756_),
    .B1(_04758_),
    .Y(_04759_));
 sky130_fd_sc_hd__or3_1 _12323_ (.A(_04750_),
    .B(_04756_),
    .C(_04758_),
    .X(_04760_));
 sky130_fd_sc_hd__nand2_1 _12324_ (.A(_04759_),
    .B(_04760_),
    .Y(_04761_));
 sky130_fd_sc_hd__a21bo_1 _12325_ (.A1(_01289_),
    .A2(_04748_),
    .B1_N(_04747_),
    .X(_04762_));
 sky130_fd_sc_hd__nand2_1 _12326_ (.A(_00460_),
    .B(_02090_),
    .Y(_04764_));
 sky130_fd_sc_hd__xnor2_2 _12327_ (.A(_04762_),
    .B(_04764_),
    .Y(_04765_));
 sky130_fd_sc_hd__and4_1 _12328_ (.A(_01066_),
    .B(_01188_),
    .C(_03414_),
    .D(_01289_),
    .X(_04766_));
 sky130_fd_sc_hd__and2b_1 _12329_ (.A_N(_04765_),
    .B(_04766_),
    .X(_04767_));
 sky130_fd_sc_hd__xnor2_1 _12330_ (.A(_04753_),
    .B(_04755_),
    .Y(_04768_));
 sky130_fd_sc_hd__nand2_1 _12331_ (.A(_04767_),
    .B(_04768_),
    .Y(_04769_));
 sky130_fd_sc_hd__o21a_1 _12332_ (.A1(_04761_),
    .A2(_04769_),
    .B1(_04759_),
    .X(_04770_));
 sky130_fd_sc_hd__xor2_1 _12333_ (.A(_04744_),
    .B(_04746_),
    .X(_04771_));
 sky130_fd_sc_hd__and2b_1 _12334_ (.A_N(_04770_),
    .B(_04771_),
    .X(_04772_));
 sky130_fd_sc_hd__a21o_1 _12335_ (.A1(_04744_),
    .A2(_04746_),
    .B1(_04772_),
    .X(_04773_));
 sky130_fd_sc_hd__xnor2_2 _12336_ (.A(_04736_),
    .B(_04773_),
    .Y(_04775_));
 sky130_fd_sc_hd__and2b_1 _12337_ (.A_N(_04771_),
    .B(_04770_),
    .X(_04776_));
 sky130_fd_sc_hd__nor2_1 _12338_ (.A(_04772_),
    .B(_04776_),
    .Y(_04777_));
 sky130_fd_sc_hd__nand4_2 _12339_ (.A(_00755_),
    .B(_01260_),
    .C(_01507_),
    .D(_01369_),
    .Y(_04778_));
 sky130_fd_sc_hd__a22o_1 _12340_ (.A1(_03762_),
    .A2(_01368_),
    .B1(_00959_),
    .B2(_03729_),
    .X(_04779_));
 sky130_fd_sc_hd__and4_1 _12341_ (.A(_03729_),
    .B(_03762_),
    .C(_01368_),
    .D(_00959_),
    .X(_04780_));
 sky130_fd_sc_hd__a31o_1 _12342_ (.A1(_01260_),
    .A2(_00605_),
    .A3(_04779_),
    .B1(_04780_),
    .X(_04781_));
 sky130_fd_sc_hd__a22o_1 _12343_ (.A1(_01260_),
    .A2(_01506_),
    .B1(_01369_),
    .B2(_00755_),
    .X(_04782_));
 sky130_fd_sc_hd__and3_1 _12344_ (.A(_04781_),
    .B(_04778_),
    .C(_04782_),
    .X(_04783_));
 sky130_fd_sc_hd__nand2_1 _12345_ (.A(_00915_),
    .B(_01664_),
    .Y(_04784_));
 sky130_fd_sc_hd__and3_1 _12346_ (.A(_00916_),
    .B(_01505_),
    .C(_04784_),
    .X(_04786_));
 sky130_fd_sc_hd__nand2_1 _12347_ (.A(_04783_),
    .B(_04786_),
    .Y(_04787_));
 sky130_fd_sc_hd__or2b_1 _12348_ (.A(_04780_),
    .B_N(_04779_),
    .X(_04788_));
 sky130_fd_sc_hd__nand2_1 _12349_ (.A(_01260_),
    .B(_00605_),
    .Y(_04789_));
 sky130_fd_sc_hd__xnor2_1 _12350_ (.A(_04788_),
    .B(_04789_),
    .Y(_04790_));
 sky130_fd_sc_hd__a22o_1 _12351_ (.A1(_03729_),
    .A2(_01506_),
    .B1(_01369_),
    .B2(_03696_),
    .X(_04791_));
 sky130_fd_sc_hd__and4_1 _12352_ (.A(_03696_),
    .B(_03729_),
    .C(_01506_),
    .D(_01369_),
    .X(_04792_));
 sky130_fd_sc_hd__a31o_1 _12353_ (.A1(_00742_),
    .A2(_00605_),
    .A3(_04791_),
    .B1(_04792_),
    .X(_04793_));
 sky130_fd_sc_hd__and2b_1 _12354_ (.A_N(_04790_),
    .B(_04793_),
    .X(_04794_));
 sky130_fd_sc_hd__a21oi_1 _12355_ (.A1(_04778_),
    .A2(_04782_),
    .B1(_04781_),
    .Y(_04795_));
 sky130_fd_sc_hd__nor2_1 _12356_ (.A(_04783_),
    .B(_04795_),
    .Y(_04797_));
 sky130_fd_sc_hd__and2_1 _12357_ (.A(_04794_),
    .B(_04797_),
    .X(_04798_));
 sky130_fd_sc_hd__and2b_1 _12358_ (.A_N(_04792_),
    .B(_04791_),
    .X(_04799_));
 sky130_fd_sc_hd__nand2_1 _12359_ (.A(_00742_),
    .B(_00605_),
    .Y(_04800_));
 sky130_fd_sc_hd__xnor2_1 _12360_ (.A(_04799_),
    .B(_04800_),
    .Y(_04801_));
 sky130_fd_sc_hd__a22o_1 _12361_ (.A1(_03729_),
    .A2(_00604_),
    .B1(_01506_),
    .B2(_03696_),
    .X(_04802_));
 sky130_fd_sc_hd__and4_1 _12362_ (.A(_03696_),
    .B(_03729_),
    .C(net46),
    .D(_01506_),
    .X(_04803_));
 sky130_fd_sc_hd__a31o_1 _12363_ (.A1(_00755_),
    .A2(_00457_),
    .A3(_04802_),
    .B1(_04803_),
    .X(_04804_));
 sky130_fd_sc_hd__nand2_1 _12364_ (.A(_00741_),
    .B(_00457_),
    .Y(_04805_));
 sky130_fd_sc_hd__xnor2_1 _12365_ (.A(_04804_),
    .B(_04805_),
    .Y(_04806_));
 sky130_fd_sc_hd__or2b_1 _12366_ (.A(_04805_),
    .B_N(_04804_),
    .X(_04808_));
 sky130_fd_sc_hd__a21bo_1 _12367_ (.A1(_04801_),
    .A2(_04806_),
    .B1_N(_04808_),
    .X(_04809_));
 sky130_fd_sc_hd__xnor2_1 _12368_ (.A(_04793_),
    .B(_04790_),
    .Y(_04810_));
 sky130_fd_sc_hd__nand2_1 _12369_ (.A(_04809_),
    .B(_04810_),
    .Y(_04811_));
 sky130_fd_sc_hd__xor2_1 _12370_ (.A(_04809_),
    .B(_04810_),
    .X(_04812_));
 sky130_fd_sc_hd__and2b_1 _12371_ (.A_N(_04803_),
    .B(_04802_),
    .X(_04813_));
 sky130_fd_sc_hd__nand2_1 _12372_ (.A(_00914_),
    .B(_00457_),
    .Y(_04814_));
 sky130_fd_sc_hd__xnor2_1 _12373_ (.A(_04813_),
    .B(_04814_),
    .Y(_04815_));
 sky130_fd_sc_hd__and4_1 _12374_ (.A(_00389_),
    .B(_00392_),
    .C(_00457_),
    .D(_00607_),
    .X(_04816_));
 sky130_fd_sc_hd__nand2_1 _12375_ (.A(_04815_),
    .B(_04816_),
    .Y(_04817_));
 sky130_fd_sc_hd__xnor2_1 _12376_ (.A(_04801_),
    .B(_04806_),
    .Y(_04819_));
 sky130_fd_sc_hd__nor2_1 _12377_ (.A(_04817_),
    .B(_04819_),
    .Y(_04820_));
 sky130_fd_sc_hd__nand2_1 _12378_ (.A(_04812_),
    .B(_04820_),
    .Y(_04821_));
 sky130_fd_sc_hd__nor2_1 _12379_ (.A(_04794_),
    .B(_04797_),
    .Y(_04822_));
 sky130_fd_sc_hd__or2_1 _12380_ (.A(_04798_),
    .B(_04822_),
    .X(_04823_));
 sky130_fd_sc_hd__a21oi_1 _12381_ (.A1(_04811_),
    .A2(_04821_),
    .B1(_04823_),
    .Y(_04824_));
 sky130_fd_sc_hd__xor2_1 _12382_ (.A(_04783_),
    .B(_04786_),
    .X(_04825_));
 sky130_fd_sc_hd__o21ai_1 _12383_ (.A1(_04798_),
    .A2(_04824_),
    .B1(_04825_),
    .Y(_04826_));
 sky130_fd_sc_hd__and3_1 _12384_ (.A(_04778_),
    .B(_04787_),
    .C(_04826_),
    .X(_04827_));
 sky130_fd_sc_hd__a22o_1 _12385_ (.A1(_00778_),
    .A2(_00571_),
    .B1(_00734_),
    .B2(_00782_),
    .X(_04828_));
 sky130_fd_sc_hd__and4_1 _12386_ (.A(_00782_),
    .B(_00613_),
    .C(_00571_),
    .D(_00734_),
    .X(_04830_));
 sky130_fd_sc_hd__a31o_1 _12387_ (.A1(_00374_),
    .A2(_01584_),
    .A3(_04828_),
    .B1(_04830_),
    .X(_04831_));
 sky130_fd_sc_hd__nand4_1 _12388_ (.A(_00784_),
    .B(_00779_),
    .C(_01586_),
    .D(_01584_),
    .Y(_04832_));
 sky130_fd_sc_hd__a22o_1 _12389_ (.A1(_00779_),
    .A2(_01586_),
    .B1(_01584_),
    .B2(_00784_),
    .X(_04833_));
 sky130_fd_sc_hd__and3_1 _12390_ (.A(_04831_),
    .B(_04832_),
    .C(_04833_),
    .X(_04834_));
 sky130_fd_sc_hd__nand2_1 _12391_ (.A(_01518_),
    .B(_01601_),
    .Y(_04835_));
 sky130_fd_sc_hd__and3_1 _12392_ (.A(_01517_),
    .B(_01780_),
    .C(_04835_),
    .X(_04836_));
 sky130_fd_sc_hd__xnor2_1 _12393_ (.A(_04834_),
    .B(_04836_),
    .Y(_04837_));
 sky130_fd_sc_hd__a22o_1 _12394_ (.A1(_00778_),
    .A2(_00413_),
    .B1(_00571_),
    .B2(_00782_),
    .X(_04838_));
 sky130_fd_sc_hd__and4_1 _12395_ (.A(_00782_),
    .B(_00613_),
    .C(_00413_),
    .D(_00571_),
    .X(_04839_));
 sky130_fd_sc_hd__a31o_1 _12396_ (.A1(_00374_),
    .A2(_01272_),
    .A3(_04838_),
    .B1(_04839_),
    .X(_04841_));
 sky130_fd_sc_hd__and2b_1 _12397_ (.A_N(_04830_),
    .B(_04828_),
    .X(_04842_));
 sky130_fd_sc_hd__nand2_1 _12398_ (.A(_00374_),
    .B(_01584_),
    .Y(_04843_));
 sky130_fd_sc_hd__xnor2_2 _12399_ (.A(_04842_),
    .B(_04843_),
    .Y(_04844_));
 sky130_fd_sc_hd__a21oi_1 _12400_ (.A1(_04832_),
    .A2(_04833_),
    .B1(_04831_),
    .Y(_04845_));
 sky130_fd_sc_hd__nor2_1 _12401_ (.A(_04834_),
    .B(_04845_),
    .Y(_04846_));
 sky130_fd_sc_hd__a21oi_1 _12402_ (.A1(_04841_),
    .A2(_04844_),
    .B1(_04846_),
    .Y(_04847_));
 sky130_fd_sc_hd__and2b_1 _12403_ (.A_N(_04839_),
    .B(_04838_),
    .X(_04848_));
 sky130_fd_sc_hd__nand2_1 _12404_ (.A(_00374_),
    .B(_01272_),
    .Y(_04849_));
 sky130_fd_sc_hd__xnor2_1 _12405_ (.A(_04848_),
    .B(_04849_),
    .Y(_04850_));
 sky130_fd_sc_hd__a22o_1 _12406_ (.A1(_00782_),
    .A2(_00413_),
    .B1(_00571_),
    .B2(_00373_),
    .X(_04852_));
 sky130_fd_sc_hd__and4_1 _12407_ (.A(_00373_),
    .B(_00782_),
    .C(_00413_),
    .D(_00571_),
    .X(_04853_));
 sky130_fd_sc_hd__a31o_1 _12408_ (.A1(_04059_),
    .A2(_01272_),
    .A3(_04852_),
    .B1(_04853_),
    .X(_04854_));
 sky130_fd_sc_hd__nand2_1 _12409_ (.A(_04059_),
    .B(_01584_),
    .Y(_04855_));
 sky130_fd_sc_hd__xnor2_1 _12410_ (.A(_04854_),
    .B(_04855_),
    .Y(_04856_));
 sky130_fd_sc_hd__and3_1 _12411_ (.A(_00378_),
    .B(_01584_),
    .C(_04854_),
    .X(_04857_));
 sky130_fd_sc_hd__a21o_1 _12412_ (.A1(_04850_),
    .A2(_04856_),
    .B1(_04857_),
    .X(_04858_));
 sky130_fd_sc_hd__xor2_1 _12413_ (.A(_04841_),
    .B(_04844_),
    .X(_04859_));
 sky130_fd_sc_hd__xnor2_1 _12414_ (.A(_04858_),
    .B(_04859_),
    .Y(_04860_));
 sky130_fd_sc_hd__or2b_2 _12415_ (.A(_04853_),
    .B_N(_04852_),
    .X(_04861_));
 sky130_fd_sc_hd__nand2_2 _12416_ (.A(_00378_),
    .B(_01586_),
    .Y(_04863_));
 sky130_fd_sc_hd__xnor2_4 _12417_ (.A(_04861_),
    .B(_04863_),
    .Y(_04864_));
 sky130_fd_sc_hd__and4_2 _12418_ (.A(_00375_),
    .B(_00378_),
    .C(_00414_),
    .D(_00572_),
    .X(_04865_));
 sky130_fd_sc_hd__and2b_1 _12419_ (.A_N(_04864_),
    .B(_04865_),
    .X(_04866_));
 sky130_fd_sc_hd__xor2_1 _12420_ (.A(_04850_),
    .B(_04856_),
    .X(_04867_));
 sky130_fd_sc_hd__nand2_1 _12421_ (.A(_04866_),
    .B(_04867_),
    .Y(_04868_));
 sky130_fd_sc_hd__nor2_1 _12422_ (.A(_04860_),
    .B(_04868_),
    .Y(_04869_));
 sky130_fd_sc_hd__a21oi_1 _12423_ (.A1(_04858_),
    .A2(_04859_),
    .B1(_04869_),
    .Y(_04870_));
 sky130_fd_sc_hd__and3_1 _12424_ (.A(_04841_),
    .B(_04844_),
    .C(_04846_),
    .X(_04871_));
 sky130_fd_sc_hd__o21ba_1 _12425_ (.A1(_04847_),
    .A2(_04870_),
    .B1_N(_04871_),
    .X(_04872_));
 sky130_fd_sc_hd__a21bo_1 _12426_ (.A1(_04834_),
    .A2(_04836_),
    .B1_N(_04832_),
    .X(_04874_));
 sky130_fd_sc_hd__o21ba_1 _12427_ (.A1(_04837_),
    .A2(_04872_),
    .B1_N(_04874_),
    .X(_04875_));
 sky130_fd_sc_hd__or2_1 _12428_ (.A(_04827_),
    .B(_04875_),
    .X(_04876_));
 sky130_fd_sc_hd__xor2_1 _12429_ (.A(_04761_),
    .B(_04769_),
    .X(_04877_));
 sky130_fd_sc_hd__and2b_1 _12430_ (.A_N(_04876_),
    .B(_04877_),
    .X(_04878_));
 sky130_fd_sc_hd__nand2_1 _12431_ (.A(_04777_),
    .B(_04878_),
    .Y(_04879_));
 sky130_fd_sc_hd__or2_1 _12432_ (.A(_04777_),
    .B(_04878_),
    .X(_04880_));
 sky130_fd_sc_hd__and2_1 _12433_ (.A(_04879_),
    .B(_04880_),
    .X(_04881_));
 sky130_fd_sc_hd__or3_1 _12434_ (.A(_04825_),
    .B(_04798_),
    .C(_04824_),
    .X(_04882_));
 sky130_fd_sc_hd__nand2_1 _12435_ (.A(_04826_),
    .B(_04882_),
    .Y(_04883_));
 sky130_fd_sc_hd__xnor2_1 _12436_ (.A(_04837_),
    .B(_04872_),
    .Y(_04885_));
 sky130_fd_sc_hd__or2_1 _12437_ (.A(_04883_),
    .B(_04885_),
    .X(_04886_));
 sky130_fd_sc_hd__xnor2_2 _12438_ (.A(_04827_),
    .B(_04875_),
    .Y(_04887_));
 sky130_fd_sc_hd__or2_1 _12439_ (.A(_04767_),
    .B(_04768_),
    .X(_04888_));
 sky130_fd_sc_hd__nand2_1 _12440_ (.A(_04769_),
    .B(_04888_),
    .Y(_04889_));
 sky130_fd_sc_hd__a21o_1 _12441_ (.A1(_04886_),
    .A2(_04887_),
    .B1(_04889_),
    .X(_04890_));
 sky130_fd_sc_hd__o21a_1 _12442_ (.A1(_04886_),
    .A2(_04887_),
    .B1(_04890_),
    .X(_04891_));
 sky130_fd_sc_hd__xnor2_1 _12443_ (.A(_04876_),
    .B(_04877_),
    .Y(_04892_));
 sky130_fd_sc_hd__and2b_1 _12444_ (.A_N(_04891_),
    .B(_04892_),
    .X(_04893_));
 sky130_fd_sc_hd__and2b_1 _12445_ (.A_N(_04892_),
    .B(_04891_),
    .X(_04894_));
 sky130_fd_sc_hd__nor2_1 _12446_ (.A(_04893_),
    .B(_04894_),
    .Y(_04896_));
 sky130_fd_sc_hd__xor2_1 _12447_ (.A(_04886_),
    .B(_04887_),
    .X(_04897_));
 sky130_fd_sc_hd__xnor2_1 _12448_ (.A(_04889_),
    .B(_04897_),
    .Y(_04898_));
 sky130_fd_sc_hd__and3_1 _12449_ (.A(_04823_),
    .B(_04811_),
    .C(_04821_),
    .X(_04899_));
 sky130_fd_sc_hd__nor2_1 _12450_ (.A(_04824_),
    .B(_04899_),
    .Y(_04900_));
 sky130_fd_sc_hd__nor2_1 _12451_ (.A(_04871_),
    .B(_04847_),
    .Y(_04901_));
 sky130_fd_sc_hd__xnor2_1 _12452_ (.A(_04901_),
    .B(_04870_),
    .Y(_04902_));
 sky130_fd_sc_hd__nand2_1 _12453_ (.A(_04900_),
    .B(_04902_),
    .Y(_04903_));
 sky130_fd_sc_hd__xnor2_1 _12454_ (.A(_04883_),
    .B(_04885_),
    .Y(_04904_));
 sky130_fd_sc_hd__nand2_1 _12455_ (.A(_04903_),
    .B(_04904_),
    .Y(_04905_));
 sky130_fd_sc_hd__xnor2_2 _12456_ (.A(_04765_),
    .B(_04766_),
    .Y(_04907_));
 sky130_fd_sc_hd__nor2_1 _12457_ (.A(_04903_),
    .B(_04904_),
    .Y(_04908_));
 sky130_fd_sc_hd__a21o_1 _12458_ (.A1(_04905_),
    .A2(_04907_),
    .B1(_04908_),
    .X(_04909_));
 sky130_fd_sc_hd__or2_1 _12459_ (.A(_04898_),
    .B(_04909_),
    .X(_04910_));
 sky130_fd_sc_hd__and2_1 _12460_ (.A(_04903_),
    .B(_04904_),
    .X(_04911_));
 sky130_fd_sc_hd__nor2_1 _12461_ (.A(_04908_),
    .B(_04911_),
    .Y(_04912_));
 sky130_fd_sc_hd__xnor2_2 _12462_ (.A(_04907_),
    .B(_04912_),
    .Y(_04913_));
 sky130_fd_sc_hd__or2_1 _12463_ (.A(_04812_),
    .B(_04820_),
    .X(_04914_));
 sky130_fd_sc_hd__and2_1 _12464_ (.A(_04821_),
    .B(_04914_),
    .X(_04915_));
 sky130_fd_sc_hd__and2_1 _12465_ (.A(_04860_),
    .B(_04868_),
    .X(_04916_));
 sky130_fd_sc_hd__nor2_1 _12466_ (.A(_04869_),
    .B(_04916_),
    .Y(_04918_));
 sky130_fd_sc_hd__nand2_1 _12467_ (.A(_04915_),
    .B(_04918_),
    .Y(_04919_));
 sky130_fd_sc_hd__xnor2_1 _12468_ (.A(_04900_),
    .B(_04902_),
    .Y(_04920_));
 sky130_fd_sc_hd__nand2_1 _12469_ (.A(_04919_),
    .B(_04920_),
    .Y(_04921_));
 sky130_fd_sc_hd__a22oi_1 _12470_ (.A1(_02008_),
    .A2(_03414_),
    .B1(_01289_),
    .B2(_04714_),
    .Y(_04922_));
 sky130_fd_sc_hd__nor2_1 _12471_ (.A(_04766_),
    .B(_04922_),
    .Y(_04923_));
 sky130_fd_sc_hd__nor2_1 _12472_ (.A(_04919_),
    .B(_04920_),
    .Y(_04924_));
 sky130_fd_sc_hd__a21oi_2 _12473_ (.A1(_04921_),
    .A2(_04923_),
    .B1(_04924_),
    .Y(_04925_));
 sky130_fd_sc_hd__xor2_2 _12474_ (.A(_04913_),
    .B(_04925_),
    .X(_04926_));
 sky130_fd_sc_hd__and2b_1 _12475_ (.A_N(_04924_),
    .B(_04921_),
    .X(_04927_));
 sky130_fd_sc_hd__xnor2_1 _12476_ (.A(_04923_),
    .B(_04927_),
    .Y(_04929_));
 sky130_fd_sc_hd__and2_1 _12477_ (.A(_04714_),
    .B(_02008_),
    .X(_04930_));
 sky130_fd_sc_hd__or2_1 _12478_ (.A(_04915_),
    .B(_04918_),
    .X(_04931_));
 sky130_fd_sc_hd__and2_1 _12479_ (.A(_04919_),
    .B(_04931_),
    .X(_04932_));
 sky130_fd_sc_hd__and2_1 _12480_ (.A(_04817_),
    .B(_04819_),
    .X(_04933_));
 sky130_fd_sc_hd__nor2_1 _12481_ (.A(_04820_),
    .B(_04933_),
    .Y(_04934_));
 sky130_fd_sc_hd__a22o_1 _12482_ (.A1(_00777_),
    .A2(_03729_),
    .B1(_03762_),
    .B2(_00612_),
    .X(_04935_));
 sky130_fd_sc_hd__and4_1 _12483_ (.A(_00612_),
    .B(_00777_),
    .C(_00423_),
    .D(_03762_),
    .X(_04936_));
 sky130_fd_sc_hd__a31o_1 _12484_ (.A1(_00374_),
    .A2(_00741_),
    .A3(_04935_),
    .B1(_04936_),
    .X(_04937_));
 sky130_fd_sc_hd__nand4_1 _12485_ (.A(_00784_),
    .B(_00779_),
    .C(_00742_),
    .D(_00741_),
    .Y(_04938_));
 sky130_fd_sc_hd__a22o_1 _12486_ (.A1(_00779_),
    .A2(_00755_),
    .B1(_00741_),
    .B2(_00783_),
    .X(_04940_));
 sky130_fd_sc_hd__and3_1 _12487_ (.A(_04937_),
    .B(_04938_),
    .C(_04940_),
    .X(_04941_));
 sky130_fd_sc_hd__nand2_1 _12488_ (.A(_01518_),
    .B(_00914_),
    .Y(_04942_));
 sky130_fd_sc_hd__and3_1 _12489_ (.A(_01517_),
    .B(_00916_),
    .C(_04942_),
    .X(_04943_));
 sky130_fd_sc_hd__xnor2_2 _12490_ (.A(_04941_),
    .B(_04943_),
    .Y(_04944_));
 sky130_fd_sc_hd__a22o_1 _12491_ (.A1(_00613_),
    .A2(_03696_),
    .B1(_03729_),
    .B2(_00612_),
    .X(_04945_));
 sky130_fd_sc_hd__and4_1 _12492_ (.A(_00780_),
    .B(_00777_),
    .C(_03685_),
    .D(_00423_),
    .X(_04946_));
 sky130_fd_sc_hd__a31o_1 _12493_ (.A1(_00374_),
    .A2(_00755_),
    .A3(_04945_),
    .B1(_04946_),
    .X(_04947_));
 sky130_fd_sc_hd__and2b_1 _12494_ (.A_N(_04936_),
    .B(_04935_),
    .X(_04948_));
 sky130_fd_sc_hd__nand2_1 _12495_ (.A(_04037_),
    .B(_03938_),
    .Y(_04949_));
 sky130_fd_sc_hd__xnor2_1 _12496_ (.A(_04948_),
    .B(_04949_),
    .Y(_04951_));
 sky130_fd_sc_hd__a21oi_1 _12497_ (.A1(_04938_),
    .A2(_04940_),
    .B1(_04937_),
    .Y(_04952_));
 sky130_fd_sc_hd__nor2_1 _12498_ (.A(_04941_),
    .B(_04952_),
    .Y(_04953_));
 sky130_fd_sc_hd__a21oi_1 _12499_ (.A1(_04947_),
    .A2(_04951_),
    .B1(_04953_),
    .Y(_04954_));
 sky130_fd_sc_hd__a22o_1 _12500_ (.A1(_00612_),
    .A2(_03696_),
    .B1(_03729_),
    .B2(_04026_),
    .X(_04955_));
 sky130_fd_sc_hd__and4_1 _12501_ (.A(_04026_),
    .B(_00780_),
    .C(_03685_),
    .D(_00423_),
    .X(_04956_));
 sky130_fd_sc_hd__a31o_1 _12502_ (.A1(_04048_),
    .A2(_03894_),
    .A3(_04955_),
    .B1(_04956_),
    .X(_04957_));
 sky130_fd_sc_hd__and3_1 _12503_ (.A(_00378_),
    .B(_00741_),
    .C(_04957_),
    .X(_04958_));
 sky130_fd_sc_hd__or2b_1 _12504_ (.A(_04946_),
    .B_N(_04945_),
    .X(_04959_));
 sky130_fd_sc_hd__nand2_1 _12505_ (.A(_04037_),
    .B(_03773_),
    .Y(_04960_));
 sky130_fd_sc_hd__xnor2_2 _12506_ (.A(_04959_),
    .B(_04960_),
    .Y(_04962_));
 sky130_fd_sc_hd__nand2_1 _12507_ (.A(_04059_),
    .B(_03938_),
    .Y(_04963_));
 sky130_fd_sc_hd__xnor2_1 _12508_ (.A(_04957_),
    .B(_04963_),
    .Y(_04964_));
 sky130_fd_sc_hd__and2b_1 _12509_ (.A_N(_04962_),
    .B(_04964_),
    .X(_04965_));
 sky130_fd_sc_hd__xor2_1 _12510_ (.A(_04947_),
    .B(_04951_),
    .X(_04966_));
 sky130_fd_sc_hd__or3_1 _12511_ (.A(_04958_),
    .B(_04965_),
    .C(_04966_),
    .X(_04967_));
 sky130_fd_sc_hd__or2b_2 _12512_ (.A(_04956_),
    .B_N(_04955_),
    .X(_04968_));
 sky130_fd_sc_hd__nand2_2 _12513_ (.A(_04059_),
    .B(_00755_),
    .Y(_04969_));
 sky130_fd_sc_hd__xnor2_4 _12514_ (.A(_04968_),
    .B(_04969_),
    .Y(_04970_));
 sky130_fd_sc_hd__and4_2 _12515_ (.A(_00374_),
    .B(_04059_),
    .C(_03707_),
    .D(_03740_),
    .X(_04971_));
 sky130_fd_sc_hd__and2b_1 _12516_ (.A_N(_04970_),
    .B(_04971_),
    .X(_04973_));
 sky130_fd_sc_hd__xnor2_1 _12517_ (.A(_04962_),
    .B(_04964_),
    .Y(_04974_));
 sky130_fd_sc_hd__and2_1 _12518_ (.A(_04973_),
    .B(_04974_),
    .X(_04975_));
 sky130_fd_sc_hd__o21a_1 _12519_ (.A1(_04958_),
    .A2(_04965_),
    .B1(_04966_),
    .X(_04976_));
 sky130_fd_sc_hd__a21oi_2 _12520_ (.A1(_04967_),
    .A2(_04975_),
    .B1(_04976_),
    .Y(_04977_));
 sky130_fd_sc_hd__nand3_1 _12521_ (.A(_04947_),
    .B(_04951_),
    .C(_04953_),
    .Y(_04978_));
 sky130_fd_sc_hd__o21ai_2 _12522_ (.A1(_04954_),
    .A2(_04977_),
    .B1(_04978_),
    .Y(_04979_));
 sky130_fd_sc_hd__and2b_1 _12523_ (.A_N(_04944_),
    .B(_04979_),
    .X(_04980_));
 sky130_fd_sc_hd__a21bo_1 _12524_ (.A1(_04941_),
    .A2(_04943_),
    .B1_N(_04938_),
    .X(_04981_));
 sky130_fd_sc_hd__or3_1 _12525_ (.A(_04934_),
    .B(_04980_),
    .C(_04981_),
    .X(_04982_));
 sky130_fd_sc_hd__o21ai_1 _12526_ (.A1(_04980_),
    .A2(_04981_),
    .B1(_04934_),
    .Y(_04984_));
 sky130_fd_sc_hd__or2_1 _12527_ (.A(_04866_),
    .B(_04867_),
    .X(_04985_));
 sky130_fd_sc_hd__nand2_1 _12528_ (.A(_04868_),
    .B(_04985_),
    .Y(_04986_));
 sky130_fd_sc_hd__nand2_1 _12529_ (.A(_04984_),
    .B(_04986_),
    .Y(_04987_));
 sky130_fd_sc_hd__and3_1 _12530_ (.A(_04932_),
    .B(_04982_),
    .C(_04987_),
    .X(_04988_));
 sky130_fd_sc_hd__a21oi_1 _12531_ (.A1(_04982_),
    .A2(_04987_),
    .B1(_04932_),
    .Y(_04989_));
 sky130_fd_sc_hd__o21bai_1 _12532_ (.A1(_04930_),
    .A2(_04988_),
    .B1_N(_04989_),
    .Y(_04990_));
 sky130_fd_sc_hd__xor2_1 _12533_ (.A(_04929_),
    .B(_04990_),
    .X(_04991_));
 sky130_fd_sc_hd__nor2_1 _12534_ (.A(_04989_),
    .B(_04988_),
    .Y(_04992_));
 sky130_fd_sc_hd__xor2_2 _12535_ (.A(_04930_),
    .B(_04992_),
    .X(_04993_));
 sky130_fd_sc_hd__nand2_1 _12536_ (.A(_04982_),
    .B(_04984_),
    .Y(_04995_));
 sky130_fd_sc_hd__xor2_1 _12537_ (.A(_04986_),
    .B(_04995_),
    .X(_04996_));
 sky130_fd_sc_hd__or2_1 _12538_ (.A(_04815_),
    .B(_04816_),
    .X(_04997_));
 sky130_fd_sc_hd__nand2_2 _12539_ (.A(_04817_),
    .B(_04997_),
    .Y(_04998_));
 sky130_fd_sc_hd__xor2_2 _12540_ (.A(_04944_),
    .B(_04979_),
    .X(_04999_));
 sky130_fd_sc_hd__xnor2_4 _12541_ (.A(_04864_),
    .B(_04865_),
    .Y(_05000_));
 sky130_fd_sc_hd__o21ba_1 _12542_ (.A1(_04998_),
    .A2(_04999_),
    .B1_N(_05000_),
    .X(_05001_));
 sky130_fd_sc_hd__a21o_1 _12543_ (.A1(_04998_),
    .A2(_04999_),
    .B1(_05001_),
    .X(_05002_));
 sky130_fd_sc_hd__or2b_1 _12544_ (.A(_04996_),
    .B_N(_05002_),
    .X(_05003_));
 sky130_fd_sc_hd__inv_2 _12545_ (.A(_04816_),
    .Y(_05004_));
 sky130_fd_sc_hd__a22o_1 _12546_ (.A1(_00393_),
    .A2(_00459_),
    .B1(_01400_),
    .B2(_00390_),
    .X(_05006_));
 sky130_fd_sc_hd__inv_2 _12547_ (.A(_04978_),
    .Y(_05007_));
 sky130_fd_sc_hd__nor2_1 _12548_ (.A(_05007_),
    .B(_04954_),
    .Y(_05008_));
 sky130_fd_sc_hd__xnor2_1 _12549_ (.A(_05008_),
    .B(net185),
    .Y(_05009_));
 sky130_fd_sc_hd__a21o_1 _12550_ (.A1(_05004_),
    .A2(_05006_),
    .B1(_05009_),
    .X(_05010_));
 sky130_fd_sc_hd__a22oi_1 _12551_ (.A1(_00376_),
    .A2(_01188_),
    .B1(_01289_),
    .B2(_00380_),
    .Y(_05011_));
 sky130_fd_sc_hd__nor2_2 _12552_ (.A(_04865_),
    .B(_05011_),
    .Y(_05012_));
 sky130_fd_sc_hd__nand3_1 _12553_ (.A(_05004_),
    .B(_05006_),
    .C(_05009_),
    .Y(_05013_));
 sky130_fd_sc_hd__a21bo_2 _12554_ (.A1(_05010_),
    .A2(_05012_),
    .B1_N(_05013_),
    .X(_05014_));
 sky130_fd_sc_hd__xor2_2 _12555_ (.A(_04998_),
    .B(_04999_),
    .X(_05015_));
 sky130_fd_sc_hd__xnor2_4 _12556_ (.A(_05000_),
    .B(_05015_),
    .Y(_05017_));
 sky130_fd_sc_hd__xor2_4 _12557_ (.A(_05014_),
    .B(_05017_),
    .X(_05018_));
 sky130_fd_sc_hd__or2b_1 _12558_ (.A(_04976_),
    .B_N(_04967_),
    .X(_05019_));
 sky130_fd_sc_hd__xnor2_2 _12559_ (.A(_05019_),
    .B(_04975_),
    .Y(_05020_));
 sky130_fd_sc_hd__a21o_1 _12560_ (.A1(_00390_),
    .A2(_04714_),
    .B1(_05020_),
    .X(_05021_));
 sky130_fd_sc_hd__and3_1 _12561_ (.A(_00390_),
    .B(_01066_),
    .C(_05020_),
    .X(_05022_));
 sky130_fd_sc_hd__a21o_1 _12562_ (.A1(_00380_),
    .A2(_02008_),
    .B1(_05022_),
    .X(_05023_));
 sky130_fd_sc_hd__nand2_2 _12563_ (.A(_05021_),
    .B(_05023_),
    .Y(_05024_));
 sky130_fd_sc_hd__nand2_1 _12564_ (.A(_05013_),
    .B(_05010_),
    .Y(_05025_));
 sky130_fd_sc_hd__xor2_2 _12565_ (.A(_05012_),
    .B(_05025_),
    .X(_05026_));
 sky130_fd_sc_hd__or2b_1 _12566_ (.A(_05017_),
    .B_N(_05014_),
    .X(_05028_));
 sky130_fd_sc_hd__o31ai_4 _12567_ (.A1(_05018_),
    .A2(_05024_),
    .A3(_05026_),
    .B1(_05028_),
    .Y(_05029_));
 sky130_fd_sc_hd__and2b_1 _12568_ (.A_N(_05002_),
    .B(_04996_),
    .X(_05030_));
 sky130_fd_sc_hd__a21o_1 _12569_ (.A1(_05003_),
    .A2(_05029_),
    .B1(_05030_),
    .X(_05031_));
 sky130_fd_sc_hd__nor2_1 _12570_ (.A(_04929_),
    .B(_04990_),
    .Y(_05032_));
 sky130_fd_sc_hd__a31o_1 _12571_ (.A1(_04991_),
    .A2(_04993_),
    .A3(_05031_),
    .B1(_05032_),
    .X(_05033_));
 sky130_fd_sc_hd__nor2_1 _12572_ (.A(_04913_),
    .B(_04925_),
    .Y(_05034_));
 sky130_fd_sc_hd__a221o_1 _12573_ (.A1(_04898_),
    .A2(_04909_),
    .B1(_04926_),
    .B2(_05033_),
    .C1(_05034_),
    .X(_05035_));
 sky130_fd_sc_hd__a31o_1 _12574_ (.A1(_04896_),
    .A2(_04910_),
    .A3(_05035_),
    .B1(_04893_),
    .X(_05036_));
 sky130_fd_sc_hd__a21boi_1 _12575_ (.A1(_04881_),
    .A2(_05036_),
    .B1_N(_04879_),
    .Y(_05037_));
 sky130_fd_sc_hd__xor2_2 _12576_ (.A(_04775_),
    .B(net155),
    .X(_05039_));
 sky130_fd_sc_hd__and4_1 _12577_ (.A(_00389_),
    .B(_00393_),
    .C(_01934_),
    .D(_02169_),
    .X(_05040_));
 sky130_fd_sc_hd__inv_2 _12578_ (.A(_05040_),
    .Y(_05041_));
 sky130_fd_sc_hd__a22o_1 _12579_ (.A1(_00393_),
    .A2(_02758_),
    .B1(_02720_),
    .B2(_00390_),
    .X(_05042_));
 sky130_fd_sc_hd__and4_1 _12580_ (.A(_03740_),
    .B(_00742_),
    .C(_02849_),
    .D(_02304_),
    .X(_05043_));
 sky130_fd_sc_hd__a22o_1 _12581_ (.A1(_00742_),
    .A2(_02849_),
    .B1(_02304_),
    .B2(_00392_),
    .X(_05044_));
 sky130_fd_sc_hd__or2b_1 _12582_ (.A(_05043_),
    .B_N(_05044_),
    .X(_05045_));
 sky130_fd_sc_hd__nand2_1 _12583_ (.A(_00745_),
    .B(_01412_),
    .Y(_05046_));
 sky130_fd_sc_hd__xnor2_1 _12584_ (.A(_05045_),
    .B(_05046_),
    .Y(_05047_));
 sky130_fd_sc_hd__a22o_1 _12585_ (.A1(_03740_),
    .A2(_02158_),
    .B1(_02304_),
    .B2(_03707_),
    .X(_05048_));
 sky130_fd_sc_hd__and4_1 _12586_ (.A(_03707_),
    .B(_03740_),
    .C(_02158_),
    .D(_02304_),
    .X(_05050_));
 sky130_fd_sc_hd__a31o_1 _12587_ (.A1(_00915_),
    .A2(_01412_),
    .A3(_05048_),
    .B1(_05050_),
    .X(_05051_));
 sky130_fd_sc_hd__or2b_1 _12588_ (.A(_05047_),
    .B_N(_05051_),
    .X(_05052_));
 sky130_fd_sc_hd__a31o_1 _12589_ (.A1(_00745_),
    .A2(_01412_),
    .A3(_05044_),
    .B1(_05043_),
    .X(_05053_));
 sky130_fd_sc_hd__nand4_2 _12590_ (.A(_00915_),
    .B(_00916_),
    .C(_02855_),
    .D(_02857_),
    .Y(_05054_));
 sky130_fd_sc_hd__a22o_1 _12591_ (.A1(_00745_),
    .A2(_02855_),
    .B1(_02857_),
    .B2(_00914_),
    .X(_05055_));
 sky130_fd_sc_hd__and3_1 _12592_ (.A(_05053_),
    .B(_05054_),
    .C(_05055_),
    .X(_05056_));
 sky130_fd_sc_hd__a21oi_1 _12593_ (.A1(_05054_),
    .A2(_05055_),
    .B1(_05053_),
    .Y(_05057_));
 sky130_fd_sc_hd__nor2_1 _12594_ (.A(_05056_),
    .B(_05057_),
    .Y(_05058_));
 sky130_fd_sc_hd__xor2_2 _12595_ (.A(_05052_),
    .B(_05058_),
    .X(_05059_));
 sky130_fd_sc_hd__nand2_1 _12596_ (.A(_00745_),
    .B(_01059_),
    .Y(_05061_));
 sky130_fd_sc_hd__a22o_1 _12597_ (.A1(_03740_),
    .A2(_01411_),
    .B1(_02849_),
    .B2(_03707_),
    .X(_05062_));
 sky130_fd_sc_hd__and4_1 _12598_ (.A(_03707_),
    .B(_03740_),
    .C(_01411_),
    .D(_02849_),
    .X(_05063_));
 sky130_fd_sc_hd__a31o_1 _12599_ (.A1(_00914_),
    .A2(_01059_),
    .A3(_05062_),
    .B1(_05063_),
    .X(_05064_));
 sky130_fd_sc_hd__or2b_1 _12600_ (.A(_05061_),
    .B_N(_05064_),
    .X(_05065_));
 sky130_fd_sc_hd__and2b_1 _12601_ (.A_N(_05050_),
    .B(_05048_),
    .X(_05066_));
 sky130_fd_sc_hd__nand2_1 _12602_ (.A(_00914_),
    .B(_01412_),
    .Y(_05067_));
 sky130_fd_sc_hd__xnor2_1 _12603_ (.A(_05066_),
    .B(_05067_),
    .Y(_05068_));
 sky130_fd_sc_hd__xnor2_1 _12604_ (.A(_05064_),
    .B(_05061_),
    .Y(_05069_));
 sky130_fd_sc_hd__nand2_1 _12605_ (.A(_05068_),
    .B(_05069_),
    .Y(_05070_));
 sky130_fd_sc_hd__xor2_1 _12606_ (.A(_05051_),
    .B(_05047_),
    .X(_05072_));
 sky130_fd_sc_hd__nand3_1 _12607_ (.A(_05065_),
    .B(_05070_),
    .C(_05072_),
    .Y(_05073_));
 sky130_fd_sc_hd__and2b_1 _12608_ (.A_N(_05063_),
    .B(_05062_),
    .X(_05074_));
 sky130_fd_sc_hd__nand2_1 _12609_ (.A(_00915_),
    .B(_01059_),
    .Y(_05075_));
 sky130_fd_sc_hd__xnor2_1 _12610_ (.A(_05074_),
    .B(_05075_),
    .Y(_05076_));
 sky130_fd_sc_hd__and4_1 _12611_ (.A(_00389_),
    .B(_00393_),
    .C(_01060_),
    .D(_01412_),
    .X(_05077_));
 sky130_fd_sc_hd__nand2_1 _12612_ (.A(_05076_),
    .B(_05077_),
    .Y(_05078_));
 sky130_fd_sc_hd__xnor2_1 _12613_ (.A(_05068_),
    .B(_05069_),
    .Y(_05079_));
 sky130_fd_sc_hd__nor2_1 _12614_ (.A(_05078_),
    .B(_05079_),
    .Y(_05080_));
 sky130_fd_sc_hd__a21oi_1 _12615_ (.A1(_05065_),
    .A2(_05070_),
    .B1(_05072_),
    .Y(_05081_));
 sky130_fd_sc_hd__a21oi_1 _12616_ (.A1(_05073_),
    .A2(_05080_),
    .B1(_05081_),
    .Y(_05083_));
 sky130_fd_sc_hd__xor2_1 _12617_ (.A(_05059_),
    .B(_05083_),
    .X(_05084_));
 sky130_fd_sc_hd__a21oi_1 _12618_ (.A1(_05041_),
    .A2(_05042_),
    .B1(_05084_),
    .Y(_05085_));
 sky130_fd_sc_hd__and4_1 _12619_ (.A(_00415_),
    .B(_00575_),
    .C(_01060_),
    .D(_01413_),
    .X(_05086_));
 sky130_fd_sc_hd__a22oi_1 _12620_ (.A1(_01289_),
    .A2(_01061_),
    .B1(_01414_),
    .B2(_01188_),
    .Y(_05087_));
 sky130_fd_sc_hd__or2_2 _12621_ (.A(_05086_),
    .B(_05087_),
    .X(_05088_));
 sky130_fd_sc_hd__and3_1 _12622_ (.A(_05041_),
    .B(_05042_),
    .C(_05084_),
    .X(_05089_));
 sky130_fd_sc_hd__o21bai_2 _12623_ (.A1(_05085_),
    .A2(_05088_),
    .B1_N(_05089_),
    .Y(_05090_));
 sky130_fd_sc_hd__and3_1 _12624_ (.A(_00414_),
    .B(_00572_),
    .C(_02849_),
    .X(_05091_));
 sky130_fd_sc_hd__a22o_1 _12625_ (.A1(_00572_),
    .A2(_01411_),
    .B1(_02306_),
    .B2(_00414_),
    .X(_05092_));
 sky130_fd_sc_hd__a21bo_1 _12626_ (.A1(_01413_),
    .A2(_05091_),
    .B1_N(_05092_),
    .X(_05094_));
 sky130_fd_sc_hd__nand2_1 _12627_ (.A(_01600_),
    .B(_01060_),
    .Y(_05095_));
 sky130_fd_sc_hd__xor2_1 _12628_ (.A(_05094_),
    .B(_05095_),
    .X(_05096_));
 sky130_fd_sc_hd__nand2_1 _12629_ (.A(_05096_),
    .B(_05086_),
    .Y(_05097_));
 sky130_fd_sc_hd__or2_1 _12630_ (.A(_05096_),
    .B(_05086_),
    .X(_05098_));
 sky130_fd_sc_hd__nand2_1 _12631_ (.A(_05097_),
    .B(_05098_),
    .Y(_05099_));
 sky130_fd_sc_hd__and3_1 _12632_ (.A(_00389_),
    .B(_00392_),
    .C(_02723_),
    .X(_05100_));
 sky130_fd_sc_hd__a22o_1 _12633_ (.A1(_00392_),
    .A2(_02168_),
    .B1(_02723_),
    .B2(_00389_),
    .X(_05101_));
 sky130_fd_sc_hd__a21bo_1 _12634_ (.A1(_02168_),
    .A2(_05100_),
    .B1_N(_05101_),
    .X(_05102_));
 sky130_fd_sc_hd__nand2_1 _12635_ (.A(_00915_),
    .B(_01933_),
    .Y(_05103_));
 sky130_fd_sc_hd__xor2_1 _12636_ (.A(_05102_),
    .B(_05103_),
    .X(_05105_));
 sky130_fd_sc_hd__nand2_1 _12637_ (.A(_05105_),
    .B(_05040_),
    .Y(_05106_));
 sky130_fd_sc_hd__or2_1 _12638_ (.A(_05105_),
    .B(_05040_),
    .X(_05107_));
 sky130_fd_sc_hd__nand2_1 _12639_ (.A(_05106_),
    .B(_05107_),
    .Y(_05108_));
 sky130_fd_sc_hd__nand2_1 _12640_ (.A(_00915_),
    .B(_02855_),
    .Y(_05109_));
 sky130_fd_sc_hd__and3_1 _12641_ (.A(_00916_),
    .B(_02857_),
    .C(_05109_),
    .X(_05110_));
 sky130_fd_sc_hd__xor2_2 _12642_ (.A(_05056_),
    .B(_05110_),
    .X(_05111_));
 sky130_fd_sc_hd__and2b_1 _12643_ (.A_N(_05052_),
    .B(_05058_),
    .X(_05112_));
 sky130_fd_sc_hd__o21bai_2 _12644_ (.A1(_05059_),
    .A2(_05083_),
    .B1_N(_05112_),
    .Y(_05113_));
 sky130_fd_sc_hd__xnor2_2 _12645_ (.A(_05111_),
    .B(_05113_),
    .Y(_05114_));
 sky130_fd_sc_hd__xor2_1 _12646_ (.A(_05108_),
    .B(_05114_),
    .X(_05116_));
 sky130_fd_sc_hd__xnor2_2 _12647_ (.A(_05099_),
    .B(_05116_),
    .Y(_05117_));
 sky130_fd_sc_hd__xor2_2 _12648_ (.A(_05090_),
    .B(_05117_),
    .X(_05118_));
 sky130_fd_sc_hd__nand2_1 _12649_ (.A(_02008_),
    .B(_01061_),
    .Y(_05119_));
 sky130_fd_sc_hd__or2b_1 _12650_ (.A(_05081_),
    .B_N(_05073_),
    .X(_05120_));
 sky130_fd_sc_hd__xnor2_1 _12651_ (.A(_05120_),
    .B(_05080_),
    .Y(_05121_));
 sky130_fd_sc_hd__and3_1 _12652_ (.A(_00390_),
    .B(_02759_),
    .C(_05121_),
    .X(_05122_));
 sky130_fd_sc_hd__inv_2 _12653_ (.A(_05122_),
    .Y(_05123_));
 sky130_fd_sc_hd__a21o_1 _12654_ (.A1(_00390_),
    .A2(_02759_),
    .B1(_05121_),
    .X(_05124_));
 sky130_fd_sc_hd__a21bo_1 _12655_ (.A1(_05119_),
    .A2(_05123_),
    .B1_N(_05124_),
    .X(_05125_));
 sky130_fd_sc_hd__or2_1 _12656_ (.A(_05089_),
    .B(_05085_),
    .X(_05127_));
 sky130_fd_sc_hd__xnor2_2 _12657_ (.A(_05088_),
    .B(_05127_),
    .Y(_05128_));
 sky130_fd_sc_hd__nor2_1 _12658_ (.A(_05125_),
    .B(_05128_),
    .Y(_05129_));
 sky130_fd_sc_hd__xor2_2 _12659_ (.A(_05118_),
    .B(_05129_),
    .X(_05130_));
 sky130_fd_sc_hd__xnor2_1 _12660_ (.A(_05039_),
    .B(_05130_),
    .Y(_05131_));
 sky130_fd_sc_hd__xnor2_1 _12661_ (.A(_04725_),
    .B(_05131_),
    .Y(_05132_));
 sky130_fd_sc_hd__xor2_2 _12662_ (.A(_04881_),
    .B(_05036_),
    .X(_05133_));
 sky130_fd_sc_hd__xor2_2 _12663_ (.A(_05125_),
    .B(_05128_),
    .X(_05134_));
 sky130_fd_sc_hd__and2_1 _12664_ (.A(_04721_),
    .B(_04723_),
    .X(_05135_));
 sky130_fd_sc_hd__or2_2 _12665_ (.A(_04724_),
    .B(_05135_),
    .X(_05136_));
 sky130_fd_sc_hd__a21boi_1 _12666_ (.A1(_05133_),
    .A2(_05134_),
    .B1_N(_05136_),
    .Y(_05138_));
 sky130_fd_sc_hd__o21ba_1 _12667_ (.A1(_05133_),
    .A2(_05134_),
    .B1_N(_05138_),
    .X(_05139_));
 sky130_fd_sc_hd__or2b_1 _12668_ (.A(_05132_),
    .B_N(_05139_),
    .X(_05140_));
 sky130_fd_sc_hd__and3_1 _12669_ (.A(_04896_),
    .B(_04910_),
    .C(_05035_),
    .X(_05141_));
 sky130_fd_sc_hd__a21oi_2 _12670_ (.A1(_04910_),
    .A2(_05035_),
    .B1(_04896_),
    .Y(_05142_));
 sky130_fd_sc_hd__nand2_1 _12671_ (.A(_05124_),
    .B(_05123_),
    .Y(_05143_));
 sky130_fd_sc_hd__xnor2_1 _12672_ (.A(_05119_),
    .B(_05143_),
    .Y(_05144_));
 sky130_fd_sc_hd__nor3_1 _12673_ (.A(_05141_),
    .B(_05142_),
    .C(_05144_),
    .Y(_05145_));
 sky130_fd_sc_hd__inv_2 _12674_ (.A(_04717_),
    .Y(_05146_));
 sky130_fd_sc_hd__o211ai_1 _12675_ (.A1(_05146_),
    .A2(_04718_),
    .B1(_00381_),
    .C1(_01958_),
    .Y(_05147_));
 sky130_fd_sc_hd__a211o_1 _12676_ (.A1(_00381_),
    .A2(_01958_),
    .B1(_05146_),
    .C1(_04718_),
    .X(_05149_));
 sky130_fd_sc_hd__nand2_2 _12677_ (.A(_05147_),
    .B(_05149_),
    .Y(_05150_));
 sky130_fd_sc_hd__xor2_1 _12678_ (.A(_05133_),
    .B(_05134_),
    .X(_05151_));
 sky130_fd_sc_hd__xnor2_1 _12679_ (.A(_05136_),
    .B(_05151_),
    .Y(_05152_));
 sky130_fd_sc_hd__o21ai_1 _12680_ (.A1(_05141_),
    .A2(_05142_),
    .B1(_05144_),
    .Y(_05153_));
 sky130_fd_sc_hd__o211a_1 _12681_ (.A1(_05145_),
    .A2(_05150_),
    .B1(_05152_),
    .C1(_05153_),
    .X(_05154_));
 sky130_fd_sc_hd__inv_2 _12682_ (.A(_05154_),
    .Y(_05155_));
 sky130_fd_sc_hd__o21a_1 _12683_ (.A1(_05141_),
    .A2(_05142_),
    .B1(_05144_),
    .X(_05156_));
 sky130_fd_sc_hd__or3_1 _12684_ (.A(_05156_),
    .B(_05145_),
    .C(_05150_),
    .X(_05157_));
 sky130_fd_sc_hd__o21ai_1 _12685_ (.A1(_05156_),
    .A2(_05145_),
    .B1(_05150_),
    .Y(_05158_));
 sky130_fd_sc_hd__and2_1 _12686_ (.A(_05078_),
    .B(_05079_),
    .X(_05160_));
 sky130_fd_sc_hd__or2_1 _12687_ (.A(_05080_),
    .B(_05160_),
    .X(_05161_));
 sky130_fd_sc_hd__a21o_1 _12688_ (.A1(_04926_),
    .A2(_05033_),
    .B1(_05034_),
    .X(_05162_));
 sky130_fd_sc_hd__nand2_1 _12689_ (.A(_04898_),
    .B(_04909_),
    .Y(_05163_));
 sky130_fd_sc_hd__and2_1 _12690_ (.A(_04910_),
    .B(_05163_),
    .X(_05164_));
 sky130_fd_sc_hd__xnor2_2 _12691_ (.A(_05162_),
    .B(_05164_),
    .Y(_05165_));
 sky130_fd_sc_hd__nor2_1 _12692_ (.A(_04692_),
    .B(_04693_),
    .Y(_05166_));
 sky130_fd_sc_hd__nor2_1 _12693_ (.A(_04694_),
    .B(_05166_),
    .Y(_05167_));
 sky130_fd_sc_hd__a21boi_1 _12694_ (.A1(_05161_),
    .A2(_05165_),
    .B1_N(_05167_),
    .Y(_05168_));
 sky130_fd_sc_hd__o21ba_1 _12695_ (.A1(_05161_),
    .A2(_05165_),
    .B1_N(_05168_),
    .X(_05169_));
 sky130_fd_sc_hd__a21oi_1 _12696_ (.A1(_05157_),
    .A2(_05158_),
    .B1(_05169_),
    .Y(_05171_));
 sky130_fd_sc_hd__xnor2_1 _12697_ (.A(_05161_),
    .B(_05165_),
    .Y(_05172_));
 sky130_fd_sc_hd__xnor2_1 _12698_ (.A(_05167_),
    .B(_05172_),
    .Y(_05173_));
 sky130_fd_sc_hd__xnor2_2 _12699_ (.A(_04926_),
    .B(_05033_),
    .Y(_05174_));
 sky130_fd_sc_hd__or2_1 _12700_ (.A(_05076_),
    .B(_05077_),
    .X(_05175_));
 sky130_fd_sc_hd__nand2_1 _12701_ (.A(_05078_),
    .B(_05175_),
    .Y(_05176_));
 sky130_fd_sc_hd__nor2_1 _12702_ (.A(_05174_),
    .B(_05176_),
    .Y(_05177_));
 sky130_fd_sc_hd__xnor2_4 _12703_ (.A(_04690_),
    .B(_04691_),
    .Y(_05178_));
 sky130_fd_sc_hd__nand2_1 _12704_ (.A(_05174_),
    .B(_05176_),
    .Y(_05179_));
 sky130_fd_sc_hd__o21a_1 _12705_ (.A1(_05177_),
    .A2(_05178_),
    .B1(_05179_),
    .X(_05180_));
 sky130_fd_sc_hd__and2_1 _12706_ (.A(_05173_),
    .B(_05180_),
    .X(_05182_));
 sky130_fd_sc_hd__inv_2 _12707_ (.A(_05077_),
    .Y(_05183_));
 sky130_fd_sc_hd__and3_1 _12708_ (.A(_04991_),
    .B(_04993_),
    .C(_05031_),
    .X(_05184_));
 sky130_fd_sc_hd__a21oi_1 _12709_ (.A1(_04993_),
    .A2(_05031_),
    .B1(_04991_),
    .Y(_05185_));
 sky130_fd_sc_hd__nor2_1 _12710_ (.A(_05184_),
    .B(_05185_),
    .Y(_05186_));
 sky130_fd_sc_hd__a22o_1 _12711_ (.A1(_00393_),
    .A2(_01062_),
    .B1(_01415_),
    .B2(_00391_),
    .X(_05187_));
 sky130_fd_sc_hd__nand2_1 _12712_ (.A(_05183_),
    .B(_05187_),
    .Y(_05188_));
 sky130_fd_sc_hd__o21ai_1 _12713_ (.A1(_05184_),
    .A2(_05185_),
    .B1(_05188_),
    .Y(_05189_));
 sky130_fd_sc_hd__a22oi_2 _12714_ (.A1(_00376_),
    .A2(_01183_),
    .B1(_01252_),
    .B2(_00380_),
    .Y(_05190_));
 sky130_fd_sc_hd__nor2_2 _12715_ (.A(_04691_),
    .B(_05190_),
    .Y(_05191_));
 sky130_fd_sc_hd__a32oi_4 _12716_ (.A1(_05183_),
    .A2(_05186_),
    .A3(_05187_),
    .B1(_05189_),
    .B2(_05191_),
    .Y(_05193_));
 sky130_fd_sc_hd__xor2_2 _12717_ (.A(_05174_),
    .B(_05176_),
    .X(_05194_));
 sky130_fd_sc_hd__xnor2_4 _12718_ (.A(_05178_),
    .B(_05194_),
    .Y(_05195_));
 sky130_fd_sc_hd__xnor2_4 _12719_ (.A(_05193_),
    .B(_05195_),
    .Y(_05196_));
 sky130_fd_sc_hd__xor2_1 _12720_ (.A(_04993_),
    .B(_05031_),
    .X(_05197_));
 sky130_fd_sc_hd__nand3_1 _12721_ (.A(_00391_),
    .B(_01108_),
    .C(_05197_),
    .Y(_05198_));
 sky130_fd_sc_hd__nand2_2 _12722_ (.A(_00380_),
    .B(_01182_),
    .Y(_05199_));
 sky130_fd_sc_hd__a21o_1 _12723_ (.A1(_00391_),
    .A2(_01062_),
    .B1(_05197_),
    .X(_05200_));
 sky130_fd_sc_hd__or2b_1 _12724_ (.A(_05199_),
    .B_N(_05200_),
    .X(_05201_));
 sky130_fd_sc_hd__and2_1 _12725_ (.A(_05198_),
    .B(_05201_),
    .X(_05202_));
 sky130_fd_sc_hd__xnor2_1 _12726_ (.A(_05186_),
    .B(_05188_),
    .Y(_05204_));
 sky130_fd_sc_hd__xnor2_2 _12727_ (.A(_05191_),
    .B(_05204_),
    .Y(_05205_));
 sky130_fd_sc_hd__or2_4 _12728_ (.A(_05202_),
    .B(_05205_),
    .X(_05206_));
 sky130_fd_sc_hd__or2_1 _12729_ (.A(_05193_),
    .B(_05195_),
    .X(_05207_));
 sky130_fd_sc_hd__o21ai_4 _12730_ (.A1(_05196_),
    .A2(_05206_),
    .B1(_05207_),
    .Y(_05208_));
 sky130_fd_sc_hd__a21o_1 _12731_ (.A1(_05157_),
    .A2(_05158_),
    .B1(_05169_),
    .X(_05209_));
 sky130_fd_sc_hd__nand3_1 _12732_ (.A(_05169_),
    .B(_05157_),
    .C(_05158_),
    .Y(_05210_));
 sky130_fd_sc_hd__or2_1 _12733_ (.A(_05173_),
    .B(_05180_),
    .X(_05211_));
 sky130_fd_sc_hd__o2111a_1 _12734_ (.A1(_05182_),
    .A2(_05208_),
    .B1(_05209_),
    .C1(_05210_),
    .D1(_05211_),
    .X(_05212_));
 sky130_fd_sc_hd__o21ai_1 _12735_ (.A1(_05145_),
    .A2(_05150_),
    .B1(_05153_),
    .Y(_05213_));
 sky130_fd_sc_hd__xnor2_1 _12736_ (.A(_05152_),
    .B(_05213_),
    .Y(_05215_));
 sky130_fd_sc_hd__o21ai_2 _12737_ (.A1(_05171_),
    .A2(_05212_),
    .B1(_05215_),
    .Y(_05216_));
 sky130_fd_sc_hd__xnor2_1 _12738_ (.A(_05132_),
    .B(_05139_),
    .Y(_05217_));
 sky130_fd_sc_hd__a21bo_1 _12739_ (.A1(_05155_),
    .A2(_05216_),
    .B1_N(_05217_),
    .X(_05218_));
 sky130_fd_sc_hd__or3b_1 _12740_ (.A(_04633_),
    .B(_04635_),
    .C_N(_04637_),
    .X(_05219_));
 sky130_fd_sc_hd__and3_1 _12741_ (.A(_00783_),
    .B(_00779_),
    .C(_02133_),
    .X(_05220_));
 sky130_fd_sc_hd__a22o_1 _12742_ (.A1(_00779_),
    .A2(_01953_),
    .B1(_02134_),
    .B2(_00784_),
    .X(_05221_));
 sky130_fd_sc_hd__a21bo_1 _12743_ (.A1(_01953_),
    .A2(_05220_),
    .B1_N(_05221_),
    .X(_05222_));
 sky130_fd_sc_hd__nand2_1 _12744_ (.A(_00375_),
    .B(_03681_),
    .Y(_05223_));
 sky130_fd_sc_hd__xor2_1 _12745_ (.A(_05222_),
    .B(_05223_),
    .X(_05224_));
 sky130_fd_sc_hd__a31o_1 _12746_ (.A1(_00378_),
    .A2(_03681_),
    .A3(_04632_),
    .B1(_04630_),
    .X(_05226_));
 sky130_fd_sc_hd__nand2_1 _12747_ (.A(_00379_),
    .B(_03678_),
    .Y(_05227_));
 sky130_fd_sc_hd__xnor2_1 _12748_ (.A(_05226_),
    .B(_05227_),
    .Y(_05228_));
 sky130_fd_sc_hd__xnor2_1 _12749_ (.A(_05224_),
    .B(_05228_),
    .Y(_05229_));
 sky130_fd_sc_hd__nor2_1 _12750_ (.A(_05219_),
    .B(_05229_),
    .Y(_05230_));
 sky130_fd_sc_hd__and2_1 _12751_ (.A(_05219_),
    .B(_05229_),
    .X(_05231_));
 sky130_fd_sc_hd__or2_1 _12752_ (.A(_05230_),
    .B(_05231_),
    .X(_05232_));
 sky130_fd_sc_hd__and3_1 _12753_ (.A(_01507_),
    .B(_01504_),
    .C(_01248_),
    .X(_05233_));
 sky130_fd_sc_hd__a22o_1 _12754_ (.A1(_01504_),
    .A2(_01179_),
    .B1(_01254_),
    .B2(_01507_),
    .X(_05234_));
 sky130_fd_sc_hd__a21bo_1 _12755_ (.A1(_01180_),
    .A2(_05233_),
    .B1_N(_05234_),
    .X(_05235_));
 sky130_fd_sc_hd__nand2_1 _12756_ (.A(_00607_),
    .B(_03738_),
    .Y(_05237_));
 sky130_fd_sc_hd__xor2_1 _12757_ (.A(_05235_),
    .B(_05237_),
    .X(_05238_));
 sky130_fd_sc_hd__a31o_1 _12758_ (.A1(_00457_),
    .A2(_03738_),
    .A3(_04640_),
    .B1(_04639_),
    .X(_05239_));
 sky130_fd_sc_hd__nand2_1 _12759_ (.A(_00457_),
    .B(_03744_),
    .Y(_05240_));
 sky130_fd_sc_hd__xnor2_1 _12760_ (.A(_05239_),
    .B(_05240_),
    .Y(_05241_));
 sky130_fd_sc_hd__xnor2_1 _12761_ (.A(_05238_),
    .B(_05241_),
    .Y(_05242_));
 sky130_fd_sc_hd__nor3_1 _12762_ (.A(_04645_),
    .B(_04646_),
    .C(_05242_),
    .Y(_05243_));
 sky130_fd_sc_hd__and2b_1 _12763_ (.A_N(_04647_),
    .B(_05242_),
    .X(_05244_));
 sky130_fd_sc_hd__or2_1 _12764_ (.A(_05243_),
    .B(_05244_),
    .X(_05245_));
 sky130_fd_sc_hd__or2b_1 _12765_ (.A(_04661_),
    .B_N(_04698_),
    .X(_05246_));
 sky130_fd_sc_hd__nand4_2 _12766_ (.A(_05245_),
    .B(_04654_),
    .C(_04659_),
    .D(_05246_),
    .Y(_05248_));
 sky130_fd_sc_hd__a31o_1 _12767_ (.A1(_04654_),
    .A2(_04659_),
    .A3(_05246_),
    .B1(_05245_),
    .X(_05249_));
 sky130_fd_sc_hd__nand2_1 _12768_ (.A(_05248_),
    .B(_05249_),
    .Y(_05250_));
 sky130_fd_sc_hd__xor2_1 _12769_ (.A(_05232_),
    .B(_05250_),
    .X(_05251_));
 sky130_fd_sc_hd__o21ba_1 _12770_ (.A1(_04649_),
    .A2(_04699_),
    .B1_N(_04638_),
    .X(_05252_));
 sky130_fd_sc_hd__a21oi_1 _12771_ (.A1(_04649_),
    .A2(_04699_),
    .B1(_05252_),
    .Y(_05253_));
 sky130_fd_sc_hd__and2_1 _12772_ (.A(_05251_),
    .B(_05253_),
    .X(_05254_));
 sky130_fd_sc_hd__or2_1 _12773_ (.A(_05251_),
    .B(_05253_),
    .X(_05255_));
 sky130_fd_sc_hd__or2b_1 _12774_ (.A(_05254_),
    .B_N(_05255_),
    .X(_05256_));
 sky130_fd_sc_hd__a21o_1 _12775_ (.A1(_04712_),
    .A2(_04724_),
    .B1(_04711_),
    .X(_05257_));
 sky130_fd_sc_hd__xor2_2 _12776_ (.A(_05256_),
    .B(_05257_),
    .X(_05259_));
 sky130_fd_sc_hd__and2_1 _12777_ (.A(_04736_),
    .B(_04773_),
    .X(_05260_));
 sky130_fd_sc_hd__nor2_1 _12778_ (.A(_04775_),
    .B(_05037_),
    .Y(_05261_));
 sky130_fd_sc_hd__a31o_1 _12779_ (.A1(_04728_),
    .A2(_04732_),
    .A3(_04735_),
    .B1(_04729_),
    .X(_05262_));
 sky130_fd_sc_hd__a22o_1 _12780_ (.A1(_00572_),
    .A2(_02849_),
    .B1(_02305_),
    .B2(_00414_),
    .X(_05263_));
 sky130_fd_sc_hd__a21bo_1 _12781_ (.A1(_02305_),
    .A2(_05091_),
    .B1_N(_05263_),
    .X(_05264_));
 sky130_fd_sc_hd__nand2_1 _12782_ (.A(_01600_),
    .B(_01412_),
    .Y(_05265_));
 sky130_fd_sc_hd__xor2_1 _12783_ (.A(_05264_),
    .B(_05265_),
    .X(_05266_));
 sky130_fd_sc_hd__and4_1 _12784_ (.A(_00414_),
    .B(_00572_),
    .C(_01411_),
    .D(_02849_),
    .X(_05267_));
 sky130_fd_sc_hd__a31o_1 _12785_ (.A1(_01586_),
    .A2(_01059_),
    .A3(_05092_),
    .B1(_05267_),
    .X(_05268_));
 sky130_fd_sc_hd__nand2_1 _12786_ (.A(_01585_),
    .B(_01059_),
    .Y(_05270_));
 sky130_fd_sc_hd__xnor2_1 _12787_ (.A(_05268_),
    .B(_05270_),
    .Y(_05271_));
 sky130_fd_sc_hd__xnor2_1 _12788_ (.A(_05266_),
    .B(_05271_),
    .Y(_05272_));
 sky130_fd_sc_hd__nor2_1 _12789_ (.A(_05097_),
    .B(_05272_),
    .Y(_05273_));
 sky130_fd_sc_hd__and2_1 _12790_ (.A(_05097_),
    .B(_05272_),
    .X(_05274_));
 sky130_fd_sc_hd__or2_1 _12791_ (.A(_05273_),
    .B(_05274_),
    .X(_05275_));
 sky130_fd_sc_hd__a22o_1 _12792_ (.A1(_00392_),
    .A2(_02723_),
    .B1(_02727_),
    .B2(_00389_),
    .X(_05276_));
 sky130_fd_sc_hd__a21bo_1 _12793_ (.A1(_02728_),
    .A2(_05100_),
    .B1_N(_05276_),
    .X(_05277_));
 sky130_fd_sc_hd__nand2_1 _12794_ (.A(_00914_),
    .B(_02168_),
    .Y(_05278_));
 sky130_fd_sc_hd__xor2_1 _12795_ (.A(_05277_),
    .B(_05278_),
    .X(_05279_));
 sky130_fd_sc_hd__and4_1 _12796_ (.A(_00389_),
    .B(_00392_),
    .C(_02168_),
    .D(_02723_),
    .X(_05281_));
 sky130_fd_sc_hd__a31o_1 _12797_ (.A1(_00914_),
    .A2(_01933_),
    .A3(_05101_),
    .B1(_05281_),
    .X(_05282_));
 sky130_fd_sc_hd__nand2_1 _12798_ (.A(_00916_),
    .B(_01933_),
    .Y(_05283_));
 sky130_fd_sc_hd__xnor2_1 _12799_ (.A(_05282_),
    .B(_05283_),
    .Y(_05284_));
 sky130_fd_sc_hd__xnor2_1 _12800_ (.A(_05279_),
    .B(_05284_),
    .Y(_05285_));
 sky130_fd_sc_hd__nor2_1 _12801_ (.A(_05106_),
    .B(_05285_),
    .Y(_05286_));
 sky130_fd_sc_hd__nand2_1 _12802_ (.A(_05106_),
    .B(_05285_),
    .Y(_05287_));
 sky130_fd_sc_hd__or2b_1 _12803_ (.A(_05286_),
    .B_N(_05287_),
    .X(_05288_));
 sky130_fd_sc_hd__nand2_1 _12804_ (.A(_05056_),
    .B(_05110_),
    .Y(_05289_));
 sky130_fd_sc_hd__nand2_1 _12805_ (.A(_05111_),
    .B(_05113_),
    .Y(_05290_));
 sky130_fd_sc_hd__nand4_2 _12806_ (.A(_05288_),
    .B(_05054_),
    .C(_05289_),
    .D(_05290_),
    .Y(_05292_));
 sky130_fd_sc_hd__a31o_1 _12807_ (.A1(_05054_),
    .A2(_05289_),
    .A3(_05290_),
    .B1(_05288_),
    .X(_05293_));
 sky130_fd_sc_hd__nand2_1 _12808_ (.A(_05292_),
    .B(_05293_),
    .Y(_05294_));
 sky130_fd_sc_hd__xor2_1 _12809_ (.A(_05275_),
    .B(_05294_),
    .X(_05295_));
 sky130_fd_sc_hd__o21a_1 _12810_ (.A1(_05108_),
    .A2(_05114_),
    .B1(_05099_),
    .X(_05296_));
 sky130_fd_sc_hd__a21o_1 _12811_ (.A1(_05108_),
    .A2(_05114_),
    .B1(_05296_),
    .X(_05297_));
 sky130_fd_sc_hd__inv_2 _12812_ (.A(_05297_),
    .Y(_05298_));
 sky130_fd_sc_hd__xnor2_1 _12813_ (.A(_05295_),
    .B(_05298_),
    .Y(_05299_));
 sky130_fd_sc_hd__and2_1 _12814_ (.A(_05090_),
    .B(_05117_),
    .X(_05300_));
 sky130_fd_sc_hd__a21o_1 _12815_ (.A1(_05118_),
    .A2(_05129_),
    .B1(_05300_),
    .X(_05301_));
 sky130_fd_sc_hd__xnor2_1 _12816_ (.A(_05299_),
    .B(_05301_),
    .Y(_05303_));
 sky130_fd_sc_hd__or4_4 _12817_ (.A(_05260_),
    .B(_05261_),
    .C(_05262_),
    .D(_05303_),
    .X(_05304_));
 sky130_fd_sc_hd__o31ai_2 _12818_ (.A1(_05260_),
    .A2(_05261_),
    .A3(_05262_),
    .B1(_05303_),
    .Y(_05305_));
 sky130_fd_sc_hd__nand2_1 _12819_ (.A(_05304_),
    .B(_05305_),
    .Y(_05306_));
 sky130_fd_sc_hd__xor2_1 _12820_ (.A(_05259_),
    .B(_05306_),
    .X(_05307_));
 sky130_fd_sc_hd__nand2_1 _12821_ (.A(_05039_),
    .B(_05130_),
    .Y(_05308_));
 sky130_fd_sc_hd__nor2_1 _12822_ (.A(_05039_),
    .B(_05130_),
    .Y(_05309_));
 sky130_fd_sc_hd__a21oi_1 _12823_ (.A1(_05308_),
    .A2(_04725_),
    .B1(_05309_),
    .Y(_05310_));
 sky130_fd_sc_hd__xnor2_1 _12824_ (.A(_05307_),
    .B(_05310_),
    .Y(_05311_));
 sky130_fd_sc_hd__a21o_1 _12825_ (.A1(_05140_),
    .A2(_05218_),
    .B1(_05311_),
    .X(_05312_));
 sky130_fd_sc_hd__nand3_1 _12826_ (.A(_05311_),
    .B(_05140_),
    .C(_05218_),
    .Y(_05314_));
 sky130_fd_sc_hd__nand2_1 _12827_ (.A(_05312_),
    .B(_05314_),
    .Y(_05315_));
 sky130_fd_sc_hd__a21oi_1 _12828_ (.A1(_04601_),
    .A2(_04628_),
    .B1(_05315_),
    .Y(_05316_));
 sky130_fd_sc_hd__inv_2 _12829_ (.A(_03675_),
    .Y(_05317_));
 sky130_fd_sc_hd__a31o_1 _12830_ (.A1(_03676_),
    .A2(_05317_),
    .A3(_02792_),
    .B1(_04600_),
    .X(_05318_));
 sky130_fd_sc_hd__nand2_1 _12831_ (.A(_05307_),
    .B(_05310_),
    .Y(_05319_));
 sky130_fd_sc_hd__nand2_1 _12832_ (.A(_05295_),
    .B(_05298_),
    .Y(_05320_));
 sky130_fd_sc_hd__or2b_1 _12833_ (.A(_05299_),
    .B_N(_05301_),
    .X(_05321_));
 sky130_fd_sc_hd__or2b_1 _12834_ (.A(_05282_),
    .B_N(_05283_),
    .X(_05322_));
 sky130_fd_sc_hd__and3_1 _12835_ (.A(_00916_),
    .B(_01933_),
    .C(_05282_),
    .X(_05323_));
 sky130_fd_sc_hd__a21o_1 _12836_ (.A1(_05279_),
    .A2(_05322_),
    .B1(_05323_),
    .X(_05325_));
 sky130_fd_sc_hd__o2bb2ai_2 _12837_ (.A1_N(_02728_),
    .A2_N(_05100_),
    .B1(_05277_),
    .B2(_05278_),
    .Y(_05326_));
 sky130_fd_sc_hd__a22oi_2 _12838_ (.A1(_00742_),
    .A2(_02724_),
    .B1(_02727_),
    .B2(_00392_),
    .Y(_05327_));
 sky130_fd_sc_hd__and4_1 _12839_ (.A(_00392_),
    .B(_00742_),
    .C(_02723_),
    .D(_02727_),
    .X(_05328_));
 sky130_fd_sc_hd__nor2_1 _12840_ (.A(_05327_),
    .B(_05328_),
    .Y(_05329_));
 sky130_fd_sc_hd__nand2_1 _12841_ (.A(_00745_),
    .B(_02168_),
    .Y(_05330_));
 sky130_fd_sc_hd__xnor2_1 _12842_ (.A(_05329_),
    .B(_05330_),
    .Y(_05331_));
 sky130_fd_sc_hd__xor2_1 _12843_ (.A(_05326_),
    .B(_05331_),
    .X(_05332_));
 sky130_fd_sc_hd__xor2_1 _12844_ (.A(_05325_),
    .B(_05332_),
    .X(_05333_));
 sky130_fd_sc_hd__or2_1 _12845_ (.A(_05286_),
    .B(_05333_),
    .X(_05334_));
 sky130_fd_sc_hd__nand2_1 _12846_ (.A(_05286_),
    .B(_05333_),
    .Y(_05336_));
 sky130_fd_sc_hd__and2_1 _12847_ (.A(_05334_),
    .B(_05336_),
    .X(_05337_));
 sky130_fd_sc_hd__or2b_1 _12848_ (.A(_05268_),
    .B_N(_05270_),
    .X(_05338_));
 sky130_fd_sc_hd__and3_1 _12849_ (.A(_01585_),
    .B(_01060_),
    .C(_05268_),
    .X(_05339_));
 sky130_fd_sc_hd__a21o_1 _12850_ (.A1(_05266_),
    .A2(_05338_),
    .B1(_05339_),
    .X(_05340_));
 sky130_fd_sc_hd__o2bb2ai_1 _12851_ (.A1_N(_02857_),
    .A2_N(_05091_),
    .B1(_05264_),
    .B2(_05265_),
    .Y(_05341_));
 sky130_fd_sc_hd__a22oi_2 _12852_ (.A1(_01586_),
    .A2(_02306_),
    .B1(_02305_),
    .B2(_00574_),
    .Y(_05342_));
 sky130_fd_sc_hd__and4_1 _12853_ (.A(_00572_),
    .B(_01586_),
    .C(_02306_),
    .D(_02305_),
    .X(_05343_));
 sky130_fd_sc_hd__nor2_1 _12854_ (.A(_05342_),
    .B(_05343_),
    .Y(_05344_));
 sky130_fd_sc_hd__nand2_1 _12855_ (.A(_01584_),
    .B(_01412_),
    .Y(_05345_));
 sky130_fd_sc_hd__xnor2_1 _12856_ (.A(_05344_),
    .B(_05345_),
    .Y(_05347_));
 sky130_fd_sc_hd__xor2_1 _12857_ (.A(_05341_),
    .B(_05347_),
    .X(_05348_));
 sky130_fd_sc_hd__xor2_1 _12858_ (.A(_05340_),
    .B(_05348_),
    .X(_05349_));
 sky130_fd_sc_hd__or2_1 _12859_ (.A(_05273_),
    .B(_05349_),
    .X(_05350_));
 sky130_fd_sc_hd__nand2_1 _12860_ (.A(_05273_),
    .B(_05349_),
    .Y(_05351_));
 sky130_fd_sc_hd__and2_1 _12861_ (.A(_05350_),
    .B(_05351_),
    .X(_05352_));
 sky130_fd_sc_hd__xor2_2 _12862_ (.A(_05337_),
    .B(_05352_),
    .X(_05353_));
 sky130_fd_sc_hd__nand2_1 _12863_ (.A(_05275_),
    .B(_05293_),
    .Y(_05354_));
 sky130_fd_sc_hd__nand2_1 _12864_ (.A(_05292_),
    .B(_05354_),
    .Y(_05355_));
 sky130_fd_sc_hd__xor2_1 _12865_ (.A(_05353_),
    .B(_05355_),
    .X(_05356_));
 sky130_fd_sc_hd__nand2_1 _12866_ (.A(_02008_),
    .B(_02765_),
    .Y(_05358_));
 sky130_fd_sc_hd__xnor2_1 _12867_ (.A(_05356_),
    .B(_05358_),
    .Y(_05359_));
 sky130_fd_sc_hd__a21o_1 _12868_ (.A1(_05320_),
    .A2(_05321_),
    .B1(_05359_),
    .X(_05360_));
 sky130_fd_sc_hd__nand3_1 _12869_ (.A(_05320_),
    .B(_05321_),
    .C(_05359_),
    .Y(_05361_));
 sky130_fd_sc_hd__nand2_1 _12870_ (.A(_05360_),
    .B(_05361_),
    .Y(_05362_));
 sky130_fd_sc_hd__a21oi_1 _12871_ (.A1(_05255_),
    .A2(_05257_),
    .B1(_05254_),
    .Y(_05363_));
 sky130_fd_sc_hd__or2b_1 _12872_ (.A(_05239_),
    .B_N(_05240_),
    .X(_05364_));
 sky130_fd_sc_hd__and3_1 _12873_ (.A(_00458_),
    .B(_03748_),
    .C(_05239_),
    .X(_05365_));
 sky130_fd_sc_hd__a21o_1 _12874_ (.A1(_05238_),
    .A2(_05364_),
    .B1(_05365_),
    .X(_05366_));
 sky130_fd_sc_hd__o2bb2ai_1 _12875_ (.A1_N(_01180_),
    .A2_N(_05233_),
    .B1(_05235_),
    .B2(_05237_),
    .Y(_05367_));
 sky130_fd_sc_hd__nand2_1 _12876_ (.A(_01504_),
    .B(_01249_),
    .Y(_05369_));
 sky130_fd_sc_hd__nand2_1 _12877_ (.A(_01507_),
    .B(_02119_),
    .Y(_05370_));
 sky130_fd_sc_hd__and4_1 _12878_ (.A(_01507_),
    .B(_01369_),
    .C(_01248_),
    .D(_02117_),
    .X(_05371_));
 sky130_fd_sc_hd__a21oi_1 _12879_ (.A1(_05369_),
    .A2(_05370_),
    .B1(_05371_),
    .Y(_05372_));
 sky130_fd_sc_hd__nand2_1 _12880_ (.A(_00605_),
    .B(_02120_),
    .Y(_05373_));
 sky130_fd_sc_hd__xnor2_1 _12881_ (.A(_05372_),
    .B(_05373_),
    .Y(_05374_));
 sky130_fd_sc_hd__xor2_1 _12882_ (.A(_05367_),
    .B(_05374_),
    .X(_05375_));
 sky130_fd_sc_hd__xor2_1 _12883_ (.A(_05366_),
    .B(_05375_),
    .X(_05376_));
 sky130_fd_sc_hd__or2_1 _12884_ (.A(_05243_),
    .B(_05376_),
    .X(_05377_));
 sky130_fd_sc_hd__nand2_1 _12885_ (.A(_05243_),
    .B(_05376_),
    .Y(_05378_));
 sky130_fd_sc_hd__and2_1 _12886_ (.A(_05377_),
    .B(_05378_),
    .X(_05380_));
 sky130_fd_sc_hd__or2b_1 _12887_ (.A(_05226_),
    .B_N(_05227_),
    .X(_05381_));
 sky130_fd_sc_hd__and3_1 _12888_ (.A(_00379_),
    .B(_03678_),
    .C(_05226_),
    .X(_05382_));
 sky130_fd_sc_hd__a21o_1 _12889_ (.A1(_05224_),
    .A2(_05381_),
    .B1(_05382_),
    .X(_05383_));
 sky130_fd_sc_hd__o2bb2ai_1 _12890_ (.A1_N(_01954_),
    .A2_N(_05220_),
    .B1(_05222_),
    .B2(_05223_),
    .Y(_05384_));
 sky130_fd_sc_hd__nand2_1 _12891_ (.A(_00779_),
    .B(_02134_),
    .Y(_05385_));
 sky130_fd_sc_hd__nand2_1 _12892_ (.A(_00784_),
    .B(_02459_),
    .Y(_05386_));
 sky130_fd_sc_hd__and4_1 _12893_ (.A(_00783_),
    .B(_00778_),
    .C(_02133_),
    .D(_02459_),
    .X(_05387_));
 sky130_fd_sc_hd__a21oi_2 _12894_ (.A1(_05385_),
    .A2(_05386_),
    .B1(_05387_),
    .Y(_05388_));
 sky130_fd_sc_hd__nand2_1 _12895_ (.A(_00375_),
    .B(_02673_),
    .Y(_05389_));
 sky130_fd_sc_hd__xnor2_1 _12896_ (.A(_05388_),
    .B(_05389_),
    .Y(_05391_));
 sky130_fd_sc_hd__xor2_1 _12897_ (.A(_05384_),
    .B(_05391_),
    .X(_05392_));
 sky130_fd_sc_hd__xor2_1 _12898_ (.A(_05383_),
    .B(_05392_),
    .X(_05393_));
 sky130_fd_sc_hd__or2_1 _12899_ (.A(_05230_),
    .B(_05393_),
    .X(_05394_));
 sky130_fd_sc_hd__nand2_1 _12900_ (.A(_05230_),
    .B(_05393_),
    .Y(_05395_));
 sky130_fd_sc_hd__and2_1 _12901_ (.A(_05394_),
    .B(_05395_),
    .X(_05396_));
 sky130_fd_sc_hd__nand2_1 _12902_ (.A(_05380_),
    .B(_05396_),
    .Y(_05397_));
 sky130_fd_sc_hd__or2_1 _12903_ (.A(_05380_),
    .B(_05396_),
    .X(_05398_));
 sky130_fd_sc_hd__and2_1 _12904_ (.A(_05397_),
    .B(_05398_),
    .X(_05399_));
 sky130_fd_sc_hd__nand2_1 _12905_ (.A(_05232_),
    .B(_05249_),
    .Y(_05400_));
 sky130_fd_sc_hd__nand2_1 _12906_ (.A(_05248_),
    .B(_05400_),
    .Y(_05402_));
 sky130_fd_sc_hd__xor2_1 _12907_ (.A(_05399_),
    .B(_05402_),
    .X(_05403_));
 sky130_fd_sc_hd__nand2_1 _12908_ (.A(_04714_),
    .B(_01957_),
    .Y(_05404_));
 sky130_fd_sc_hd__xnor2_1 _12909_ (.A(_05403_),
    .B(_05404_),
    .Y(_05405_));
 sky130_fd_sc_hd__nor2_1 _12910_ (.A(_05363_),
    .B(_05405_),
    .Y(_05406_));
 sky130_fd_sc_hd__and2_1 _12911_ (.A(_05363_),
    .B(_05405_),
    .X(_05407_));
 sky130_fd_sc_hd__nor2_1 _12912_ (.A(_05406_),
    .B(_05407_),
    .Y(_05408_));
 sky130_fd_sc_hd__xnor2_1 _12913_ (.A(_05362_),
    .B(_05408_),
    .Y(_05409_));
 sky130_fd_sc_hd__nand2_1 _12914_ (.A(_05259_),
    .B(_05305_),
    .Y(_05410_));
 sky130_fd_sc_hd__and3_1 _12915_ (.A(_05409_),
    .B(_05304_),
    .C(_05410_),
    .X(_05411_));
 sky130_fd_sc_hd__a21o_1 _12916_ (.A1(_05304_),
    .A2(_05410_),
    .B1(_05409_),
    .X(_05413_));
 sky130_fd_sc_hd__or2b_1 _12917_ (.A(_05411_),
    .B_N(_05413_),
    .X(_05414_));
 sky130_fd_sc_hd__nand2_1 _12918_ (.A(_01108_),
    .B(_01183_),
    .Y(_05415_));
 sky130_fd_sc_hd__xnor2_2 _12919_ (.A(_05414_),
    .B(_05415_),
    .Y(_05416_));
 sky130_fd_sc_hd__a21oi_4 _12920_ (.A1(_05319_),
    .A2(_05312_),
    .B1(_05416_),
    .Y(_05417_));
 sky130_fd_sc_hd__and3_1 _12921_ (.A(_05416_),
    .B(_05319_),
    .C(_05312_),
    .X(_05418_));
 sky130_fd_sc_hd__nor2_1 _12922_ (.A(_05417_),
    .B(_05418_),
    .Y(_05419_));
 sky130_fd_sc_hd__xnor2_1 _12923_ (.A(_05318_),
    .B(_05419_),
    .Y(_05420_));
 sky130_fd_sc_hd__o21a_1 _12924_ (.A1(_04629_),
    .A2(_05316_),
    .B1(_05420_),
    .X(_05421_));
 sky130_fd_sc_hd__or3_1 _12925_ (.A(_05420_),
    .B(_04629_),
    .C(_05316_),
    .X(_05422_));
 sky130_fd_sc_hd__nand2b_2 _12926_ (.A_N(_05421_),
    .B(_05422_),
    .Y(_05424_));
 sky130_fd_sc_hd__nand2_1 _12927_ (.A(_04617_),
    .B(_04610_),
    .Y(_05425_));
 sky130_fd_sc_hd__xnor2_2 _12928_ (.A(_03613_),
    .B(_05425_),
    .Y(_05426_));
 sky130_fd_sc_hd__o21ai_1 _12929_ (.A1(_04575_),
    .A2(_04580_),
    .B1(_04585_),
    .Y(_05427_));
 sky130_fd_sc_hd__nand2_2 _12930_ (.A(_04491_),
    .B(_05427_),
    .Y(_05428_));
 sky130_fd_sc_hd__xnor2_4 _12931_ (.A(_04536_),
    .B(_05428_),
    .Y(_05429_));
 sky130_fd_sc_hd__xor2_2 _12932_ (.A(_05426_),
    .B(_05429_),
    .X(_05430_));
 sky130_fd_sc_hd__and3_2 _12933_ (.A(_03585_),
    .B(_03588_),
    .C(_03590_),
    .X(_05431_));
 sky130_fd_sc_hd__o21ai_1 _12934_ (.A1(_05431_),
    .A2(_03612_),
    .B1(_03619_),
    .Y(_05432_));
 sky130_fd_sc_hd__xor2_2 _12935_ (.A(_03614_),
    .B(_05432_),
    .X(_05433_));
 sky130_fd_sc_hd__inv_2 _12936_ (.A(_05433_),
    .Y(_05435_));
 sky130_fd_sc_hd__a21oi_2 _12937_ (.A1(_04566_),
    .A2(_04582_),
    .B1(_04484_),
    .Y(_05436_));
 sky130_fd_sc_hd__a2111o_1 _12938_ (.A1(_04570_),
    .A2(_04571_),
    .B1(_02473_),
    .C1(_02475_),
    .D1(_02699_),
    .X(_05437_));
 sky130_fd_sc_hd__or3_1 _12939_ (.A(_04566_),
    .B(_04583_),
    .C(_04574_),
    .X(_05438_));
 sky130_fd_sc_hd__a21o_1 _12940_ (.A1(_04573_),
    .A2(_05437_),
    .B1(_05438_),
    .X(_05439_));
 sky130_fd_sc_hd__a21o_1 _12941_ (.A1(_04570_),
    .A2(_04571_),
    .B1(_02699_),
    .X(_05440_));
 sky130_fd_sc_hd__a2111o_2 _12942_ (.A1(_02391_),
    .A2(_02150_),
    .B1(_02479_),
    .C1(_05440_),
    .D1(_05438_),
    .X(_05441_));
 sky130_fd_sc_hd__and3_2 _12943_ (.A(_05436_),
    .B(_05439_),
    .C(_05441_),
    .X(_05442_));
 sky130_fd_sc_hd__nand2_1 _12944_ (.A(_04581_),
    .B(_04403_),
    .Y(_05443_));
 sky130_fd_sc_hd__o21bai_1 _12945_ (.A1(_04402_),
    .A2(_04471_),
    .B1_N(_04401_),
    .Y(_05444_));
 sky130_fd_sc_hd__o21ai_2 _12946_ (.A1(_05442_),
    .A2(_05443_),
    .B1(_05444_),
    .Y(_05446_));
 sky130_fd_sc_hd__xnor2_4 _12947_ (.A(_05446_),
    .B(_04454_),
    .Y(_05447_));
 sky130_fd_sc_hd__nor2_1 _12948_ (.A(_05435_),
    .B(_05447_),
    .Y(_05448_));
 sky130_fd_sc_hd__or2_1 _12949_ (.A(_05430_),
    .B(_05448_),
    .X(_05449_));
 sky130_fd_sc_hd__nor2_2 _12950_ (.A(_05024_),
    .B(_05026_),
    .Y(_05450_));
 sky130_fd_sc_hd__xnor2_4 _12951_ (.A(_05018_),
    .B(_05450_),
    .Y(_05451_));
 sky130_fd_sc_hd__and2_1 _12952_ (.A(_05430_),
    .B(_05448_),
    .X(_05452_));
 sky130_fd_sc_hd__a21o_2 _12953_ (.A1(_05449_),
    .A2(_05451_),
    .B1(_05452_),
    .X(_05453_));
 sky130_fd_sc_hd__or2b_2 _12954_ (.A(_05030_),
    .B_N(_05003_),
    .X(_05454_));
 sky130_fd_sc_hd__xnor2_4 _12955_ (.A(_05454_),
    .B(_05029_),
    .Y(_05455_));
 sky130_fd_sc_hd__nor2_1 _12956_ (.A(_05426_),
    .B(_05429_),
    .Y(_05457_));
 sky130_fd_sc_hd__or2_1 _12957_ (.A(_04534_),
    .B(_04535_),
    .X(_05458_));
 sky130_fd_sc_hd__o21a_1 _12958_ (.A1(_04589_),
    .A2(_04487_),
    .B1(_05458_),
    .X(_05459_));
 sky130_fd_sc_hd__nand2_1 _12959_ (.A(_04536_),
    .B(_04454_),
    .Y(_05460_));
 sky130_fd_sc_hd__a311oi_4 _12960_ (.A1(_05436_),
    .A2(_05439_),
    .A3(_05441_),
    .B1(_05443_),
    .C1(_05460_),
    .Y(_05461_));
 sky130_fd_sc_hd__nor2_1 _12961_ (.A(_05444_),
    .B(_05460_),
    .Y(_05462_));
 sky130_fd_sc_hd__or3_4 _12962_ (.A(_05459_),
    .B(_05461_),
    .C(_05462_),
    .X(_05463_));
 sky130_fd_sc_hd__xor2_4 _12963_ (.A(_04531_),
    .B(_05463_),
    .X(_05464_));
 sky130_fd_sc_hd__or3_2 _12964_ (.A(_03536_),
    .B(_03616_),
    .C(_03621_),
    .X(_05465_));
 sky130_fd_sc_hd__xor2_2 _12965_ (.A(_05465_),
    .B(_03623_),
    .X(_05466_));
 sky130_fd_sc_hd__xnor2_1 _12966_ (.A(_05464_),
    .B(_05466_),
    .Y(_05468_));
 sky130_fd_sc_hd__inv_2 _12967_ (.A(_05468_),
    .Y(_05469_));
 sky130_fd_sc_hd__xnor2_2 _12968_ (.A(_05457_),
    .B(_05469_),
    .Y(_05470_));
 sky130_fd_sc_hd__xnor2_4 _12969_ (.A(_05455_),
    .B(_05470_),
    .Y(_05471_));
 sky130_fd_sc_hd__xor2_4 _12970_ (.A(_05453_),
    .B(_05471_),
    .X(_05472_));
 sky130_fd_sc_hd__xor2_2 _12971_ (.A(_05430_),
    .B(_05448_),
    .X(_05473_));
 sky130_fd_sc_hd__xnor2_4 _12972_ (.A(_05451_),
    .B(_05473_),
    .Y(_05474_));
 sky130_fd_sc_hd__xor2_2 _12973_ (.A(_05433_),
    .B(_05447_),
    .X(_05475_));
 sky130_fd_sc_hd__inv_2 _12974_ (.A(_05475_),
    .Y(_05476_));
 sky130_fd_sc_hd__or2_1 _12975_ (.A(_04602_),
    .B(_04607_),
    .X(_05477_));
 sky130_fd_sc_hd__o211a_1 _12976_ (.A1(_04606_),
    .A2(_04607_),
    .B1(_05477_),
    .C1(_04614_),
    .X(_05479_));
 sky130_fd_sc_hd__xor2_2 _12977_ (.A(_03602_),
    .B(_05479_),
    .X(_05480_));
 sky130_fd_sc_hd__and3_1 _12978_ (.A(_04581_),
    .B(_04584_),
    .C(_04575_),
    .X(_05481_));
 sky130_fd_sc_hd__a311oi_4 _12979_ (.A1(_04581_),
    .A2(_04584_),
    .A3(_04580_),
    .B1(_04486_),
    .C1(_05481_),
    .Y(_05482_));
 sky130_fd_sc_hd__xor2_4 _12980_ (.A(_04403_),
    .B(_05482_),
    .X(_05483_));
 sky130_fd_sc_hd__nor2_1 _12981_ (.A(_05480_),
    .B(_05483_),
    .Y(_05484_));
 sky130_fd_sc_hd__and2_1 _12982_ (.A(_05476_),
    .B(_05484_),
    .X(_05485_));
 sky130_fd_sc_hd__and2_1 _12983_ (.A(_05024_),
    .B(_05026_),
    .X(_05486_));
 sky130_fd_sc_hd__nor2_2 _12984_ (.A(_05450_),
    .B(_05486_),
    .Y(_05487_));
 sky130_fd_sc_hd__or2_1 _12985_ (.A(_05476_),
    .B(_05484_),
    .X(_05488_));
 sky130_fd_sc_hd__o21ai_4 _12986_ (.A1(_05485_),
    .A2(_05487_),
    .B1(_05488_),
    .Y(_05490_));
 sky130_fd_sc_hd__xor2_1 _12987_ (.A(_05474_),
    .B(_05490_),
    .X(_05491_));
 sky130_fd_sc_hd__and2_1 _12988_ (.A(_05472_),
    .B(_05491_),
    .X(_05492_));
 sky130_fd_sc_hd__xnor2_4 _12989_ (.A(_05431_),
    .B(_03611_),
    .Y(_05493_));
 sky130_fd_sc_hd__xnor2_4 _12990_ (.A(_04581_),
    .B(_05442_),
    .Y(_05494_));
 sky130_fd_sc_hd__xor2_2 _12991_ (.A(_05480_),
    .B(_05483_),
    .X(_05495_));
 sky130_fd_sc_hd__a21o_1 _12992_ (.A1(_05493_),
    .A2(_05494_),
    .B1(_05495_),
    .X(_05496_));
 sky130_fd_sc_hd__inv_2 _12993_ (.A(_05021_),
    .Y(_05497_));
 sky130_fd_sc_hd__o211ai_2 _12994_ (.A1(_05497_),
    .A2(_05022_),
    .B1(_00381_),
    .C1(_02008_),
    .Y(_05498_));
 sky130_fd_sc_hd__a211o_1 _12995_ (.A1(_00381_),
    .A2(_02008_),
    .B1(_05497_),
    .C1(_05022_),
    .X(_05499_));
 sky130_fd_sc_hd__nand2_4 _12996_ (.A(_05498_),
    .B(_05499_),
    .Y(_05501_));
 sky130_fd_sc_hd__a31o_1 _12997_ (.A1(_05493_),
    .A2(_05494_),
    .A3(_05495_),
    .B1(_05501_),
    .X(_05502_));
 sky130_fd_sc_hd__xnor2_1 _12998_ (.A(_05475_),
    .B(_05484_),
    .Y(_05503_));
 sky130_fd_sc_hd__xnor2_1 _12999_ (.A(_05487_),
    .B(_05503_),
    .Y(_05504_));
 sky130_fd_sc_hd__a21boi_2 _13000_ (.A1(_05496_),
    .A2(_05502_),
    .B1_N(_05504_),
    .Y(_05505_));
 sky130_fd_sc_hd__nand3b_2 _13001_ (.A_N(_05504_),
    .B(_05496_),
    .C(_05502_),
    .Y(_05506_));
 sky130_fd_sc_hd__and2b_1 _13002_ (.A_N(_05505_),
    .B(_05506_),
    .X(_05507_));
 sky130_fd_sc_hd__nor2_1 _13003_ (.A(_04973_),
    .B(_04974_),
    .Y(_05508_));
 sky130_fd_sc_hd__or2_2 _13004_ (.A(_04975_),
    .B(_05508_),
    .X(_05509_));
 sky130_fd_sc_hd__xor2_2 _13005_ (.A(_05493_),
    .B(_05494_),
    .X(_05510_));
 sky130_fd_sc_hd__a21o_1 _13006_ (.A1(_04602_),
    .A2(_04606_),
    .B1(_03578_),
    .X(_05512_));
 sky130_fd_sc_hd__o21ai_4 _13007_ (.A1(_04575_),
    .A2(_04580_),
    .B1(_04584_),
    .Y(_05513_));
 sky130_fd_sc_hd__nand3_1 _13008_ (.A(_03578_),
    .B(_04602_),
    .C(_04606_),
    .Y(_05514_));
 sky130_fd_sc_hd__or3_4 _13009_ (.A(_04584_),
    .B(_04575_),
    .C(_04580_),
    .X(_05515_));
 sky130_fd_sc_hd__and4_1 _13010_ (.A(_05512_),
    .B(_05513_),
    .C(_05514_),
    .D(_05515_),
    .X(_05516_));
 sky130_fd_sc_hd__nor2_1 _13011_ (.A(_05510_),
    .B(_05516_),
    .Y(_05517_));
 sky130_fd_sc_hd__nand2_1 _13012_ (.A(_05510_),
    .B(_05516_),
    .Y(_05518_));
 sky130_fd_sc_hd__o21a_2 _13013_ (.A1(_05509_),
    .A2(_05517_),
    .B1(_05518_),
    .X(_05519_));
 sky130_fd_sc_hd__nand2_1 _13014_ (.A(_05493_),
    .B(_05494_),
    .Y(_05520_));
 sky130_fd_sc_hd__xnor2_2 _13015_ (.A(_05520_),
    .B(_05495_),
    .Y(_05521_));
 sky130_fd_sc_hd__xnor2_4 _13016_ (.A(_05501_),
    .B(_05521_),
    .Y(_05523_));
 sky130_fd_sc_hd__xor2_4 _13017_ (.A(_05519_),
    .B(_05523_),
    .X(_05524_));
 sky130_fd_sc_hd__and3_1 _13018_ (.A(_05492_),
    .B(_05507_),
    .C(_05524_),
    .X(_05525_));
 sky130_fd_sc_hd__and2_1 _13019_ (.A(_01639_),
    .B(_02046_),
    .X(_05526_));
 sky130_fd_sc_hd__and4_1 _13020_ (.A(_01637_),
    .B(net131),
    .C(_01433_),
    .D(_02046_),
    .X(_05527_));
 sky130_fd_sc_hd__o31ai_4 _13021_ (.A1(_02049_),
    .A2(_05526_),
    .A3(_05527_),
    .B1(_02492_),
    .Y(_05528_));
 sky130_fd_sc_hd__xnor2_1 _13022_ (.A(_05510_),
    .B(_05516_),
    .Y(_05529_));
 sky130_fd_sc_hd__xnor2_1 _13023_ (.A(_05509_),
    .B(_05529_),
    .Y(_05530_));
 sky130_fd_sc_hd__a22o_1 _13024_ (.A1(_05512_),
    .A2(_05514_),
    .B1(_05515_),
    .B2(_05513_),
    .X(_05531_));
 sky130_fd_sc_hd__or2b_2 _13025_ (.A(_05516_),
    .B_N(_05531_),
    .X(_05532_));
 sky130_fd_sc_hd__nand2_1 _13026_ (.A(_04573_),
    .B(_05437_),
    .Y(_05534_));
 sky130_fd_sc_hd__a31o_1 _13027_ (.A1(_02480_),
    .A2(_04577_),
    .A3(_04579_),
    .B1(_05534_),
    .X(_05535_));
 sky130_fd_sc_hd__xnor2_4 _13028_ (.A(_04578_),
    .B(_05535_),
    .Y(_05536_));
 sky130_fd_sc_hd__o21ai_2 _13029_ (.A1(_02589_),
    .A2(_04604_),
    .B1(_03551_),
    .Y(_05537_));
 sky130_fd_sc_hd__xor2_2 _13030_ (.A(_04603_),
    .B(_05537_),
    .X(_05538_));
 sky130_fd_sc_hd__or2_2 _13031_ (.A(_05536_),
    .B(_05538_),
    .X(_05539_));
 sky130_fd_sc_hd__or2_1 _13032_ (.A(_05532_),
    .B(_05539_),
    .X(_05540_));
 sky130_fd_sc_hd__xor2_4 _13033_ (.A(_04970_),
    .B(_04971_),
    .X(_05541_));
 sky130_fd_sc_hd__a21o_1 _13034_ (.A1(_05532_),
    .A2(_05539_),
    .B1(_05541_),
    .X(_05542_));
 sky130_fd_sc_hd__and3_1 _13035_ (.A(_05530_),
    .B(_05540_),
    .C(_05542_),
    .X(_05543_));
 sky130_fd_sc_hd__a21o_1 _13036_ (.A1(_05540_),
    .A2(_05542_),
    .B1(_05530_),
    .X(_05545_));
 sky130_fd_sc_hd__and2b_2 _13037_ (.A_N(_05543_),
    .B(_05545_),
    .X(_05546_));
 sky130_fd_sc_hd__xnor2_4 _13038_ (.A(_05532_),
    .B(_05539_),
    .Y(_05547_));
 sky130_fd_sc_hd__xnor2_4 _13039_ (.A(_05541_),
    .B(_05547_),
    .Y(_05548_));
 sky130_fd_sc_hd__xor2_2 _13040_ (.A(_05536_),
    .B(_05538_),
    .X(_05549_));
 sky130_fd_sc_hd__inv_2 _13041_ (.A(_04604_),
    .Y(_05550_));
 sky130_fd_sc_hd__mux2_1 _13042_ (.A0(_05550_),
    .A1(_04605_),
    .S(_02589_),
    .X(_05551_));
 sky130_fd_sc_hd__or2b_1 _13043_ (.A(_04579_),
    .B_N(_04572_),
    .X(_05552_));
 sky130_fd_sc_hd__nand2_1 _13044_ (.A(_04573_),
    .B(_05552_),
    .Y(_05553_));
 sky130_fd_sc_hd__mux2_4 _13045_ (.A0(_04579_),
    .A1(_05553_),
    .S(_02701_),
    .X(_05554_));
 sky130_fd_sc_hd__nor2_1 _13046_ (.A(_05551_),
    .B(_05554_),
    .Y(_05556_));
 sky130_fd_sc_hd__nand2_1 _13047_ (.A(_05549_),
    .B(_05556_),
    .Y(_05557_));
 sky130_fd_sc_hd__a22oi_2 _13048_ (.A1(_00376_),
    .A2(_00391_),
    .B1(_00393_),
    .B2(_00381_),
    .Y(_05558_));
 sky130_fd_sc_hd__nor2_4 _13049_ (.A(_04971_),
    .B(_05558_),
    .Y(_05559_));
 sky130_fd_sc_hd__o21ai_1 _13050_ (.A1(_05549_),
    .A2(_05556_),
    .B1(_05559_),
    .Y(_05560_));
 sky130_fd_sc_hd__nand2_2 _13051_ (.A(_05557_),
    .B(_05560_),
    .Y(_05561_));
 sky130_fd_sc_hd__xnor2_4 _13052_ (.A(_05548_),
    .B(_05561_),
    .Y(_05562_));
 sky130_fd_sc_hd__and2_2 _13053_ (.A(_05546_),
    .B(_05562_),
    .X(_05563_));
 sky130_fd_sc_hd__and2_1 _13054_ (.A(_05551_),
    .B(_05554_),
    .X(_05564_));
 sky130_fd_sc_hd__nor2_1 _13055_ (.A(_05556_),
    .B(_05564_),
    .Y(_05565_));
 sky130_fd_sc_hd__a21boi_2 _13056_ (.A1(_02592_),
    .A2(_02703_),
    .B1_N(_02593_),
    .Y(_05567_));
 sky130_fd_sc_hd__or2_1 _13057_ (.A(_05565_),
    .B(_05567_),
    .X(_05568_));
 sky130_fd_sc_hd__nand2_2 _13058_ (.A(_00381_),
    .B(_00391_),
    .Y(_05569_));
 sky130_fd_sc_hd__a21bo_1 _13059_ (.A1(_05565_),
    .A2(_05567_),
    .B1_N(_05569_),
    .X(_05570_));
 sky130_fd_sc_hd__xnor2_1 _13060_ (.A(_05549_),
    .B(_05556_),
    .Y(_05571_));
 sky130_fd_sc_hd__xnor2_2 _13061_ (.A(_05559_),
    .B(_05571_),
    .Y(_05572_));
 sky130_fd_sc_hd__a21oi_2 _13062_ (.A1(_05568_),
    .A2(_05570_),
    .B1(_05572_),
    .Y(_05573_));
 sky130_fd_sc_hd__and3_1 _13063_ (.A(_05572_),
    .B(_05568_),
    .C(_05570_),
    .X(_05574_));
 sky130_fd_sc_hd__nor2_2 _13064_ (.A(_05573_),
    .B(_05574_),
    .Y(_05575_));
 sky130_fd_sc_hd__xor2_2 _13065_ (.A(_05565_),
    .B(_05567_),
    .X(_05576_));
 sky130_fd_sc_hd__xnor2_4 _13066_ (.A(_05569_),
    .B(_05576_),
    .Y(_05578_));
 sky130_fd_sc_hd__xnor2_4 _13067_ (.A(_02709_),
    .B(_05578_),
    .Y(_05579_));
 sky130_fd_sc_hd__and2_1 _13068_ (.A(_05575_),
    .B(_05579_),
    .X(_05580_));
 sky130_fd_sc_hd__nand2_1 _13069_ (.A(_05563_),
    .B(_05580_),
    .Y(_05581_));
 sky130_fd_sc_hd__nand2_1 _13070_ (.A(_02491_),
    .B(_02713_),
    .Y(_05582_));
 sky130_fd_sc_hd__a211o_1 _13071_ (.A1(_02483_),
    .A2(_02484_),
    .B1(_02485_),
    .C1(_02486_),
    .X(_05583_));
 sky130_fd_sc_hd__o31ai_1 _13072_ (.A1(_02055_),
    .A2(_02272_),
    .A3(_02488_),
    .B1(_05583_),
    .Y(_05584_));
 sky130_fd_sc_hd__and3_1 _13073_ (.A(_02709_),
    .B(_02710_),
    .C(_05584_),
    .X(_05585_));
 sky130_fd_sc_hd__a41o_1 _13074_ (.A1(_02273_),
    .A2(_02491_),
    .A3(_02493_),
    .A4(_02713_),
    .B1(_05585_),
    .X(_05586_));
 sky130_fd_sc_hd__nand3_1 _13075_ (.A(_05563_),
    .B(_05580_),
    .C(_05586_),
    .Y(_05587_));
 sky130_fd_sc_hd__inv_2 _13076_ (.A(_05573_),
    .Y(_05589_));
 sky130_fd_sc_hd__a21oi_1 _13077_ (.A1(_02704_),
    .A2(_02705_),
    .B1(_02707_),
    .Y(_05590_));
 sky130_fd_sc_hd__a21o_1 _13078_ (.A1(_05590_),
    .A2(_05578_),
    .B1(_05574_),
    .X(_05591_));
 sky130_fd_sc_hd__or2b_2 _13079_ (.A(_05548_),
    .B_N(_05561_),
    .X(_05592_));
 sky130_fd_sc_hd__a21oi_2 _13080_ (.A1(_05545_),
    .A2(_05592_),
    .B1(_05543_),
    .Y(_05593_));
 sky130_fd_sc_hd__a31oi_2 _13081_ (.A1(_05563_),
    .A2(_05589_),
    .A3(_05591_),
    .B1(_05593_),
    .Y(_05594_));
 sky130_fd_sc_hd__o311ai_4 _13082_ (.A1(_05528_),
    .A2(_05581_),
    .A3(_05582_),
    .B1(_05587_),
    .C1(_05594_),
    .Y(_05595_));
 sky130_fd_sc_hd__or2_1 _13083_ (.A(_05519_),
    .B(_05523_),
    .X(_05596_));
 sky130_fd_sc_hd__a21oi_2 _13084_ (.A1(_05506_),
    .A2(_05596_),
    .B1(_05505_),
    .Y(_05597_));
 sky130_fd_sc_hd__nand2_1 _13085_ (.A(_05453_),
    .B(_05471_),
    .Y(_05598_));
 sky130_fd_sc_hd__or2_1 _13086_ (.A(_05474_),
    .B(_05490_),
    .X(_05600_));
 sky130_fd_sc_hd__nor2_1 _13087_ (.A(_05453_),
    .B(_05471_),
    .Y(_05601_));
 sky130_fd_sc_hd__a21o_1 _13088_ (.A1(_05598_),
    .A2(_05600_),
    .B1(_05601_),
    .X(_05602_));
 sky130_fd_sc_hd__a21bo_1 _13089_ (.A1(_05492_),
    .A2(_05597_),
    .B1_N(_05602_),
    .X(_05603_));
 sky130_fd_sc_hd__a21oi_1 _13090_ (.A1(_05525_),
    .A2(_05595_),
    .B1(_05603_),
    .Y(_05604_));
 sky130_fd_sc_hd__xnor2_2 _13091_ (.A(_04626_),
    .B(_04627_),
    .Y(_05605_));
 sky130_fd_sc_hd__inv_2 _13092_ (.A(_03672_),
    .Y(_05606_));
 sky130_fd_sc_hd__o31a_1 _13093_ (.A1(_03456_),
    .A2(_03496_),
    .A3(_03625_),
    .B1(_05606_),
    .X(_05607_));
 sky130_fd_sc_hd__xnor2_2 _13094_ (.A(_03668_),
    .B(_05607_),
    .Y(_05608_));
 sky130_fd_sc_hd__nor3b_1 _13095_ (.A(_03956_),
    .B(_04025_),
    .C_N(_04545_),
    .Y(_05609_));
 sky130_fd_sc_hd__nand2_1 _13096_ (.A(_04548_),
    .B(_04550_),
    .Y(_05611_));
 sky130_fd_sc_hd__o21a_1 _13097_ (.A1(_04592_),
    .A2(_04588_),
    .B1(_05611_),
    .X(_05612_));
 sky130_fd_sc_hd__or2_1 _13098_ (.A(_04025_),
    .B(_04546_),
    .X(_05613_));
 sky130_fd_sc_hd__inv_2 _13099_ (.A(_05613_),
    .Y(_05614_));
 sky130_fd_sc_hd__and2_1 _13100_ (.A(_05612_),
    .B(_05614_),
    .X(_05615_));
 sky130_fd_sc_hd__and2_1 _13101_ (.A(_04551_),
    .B(_04531_),
    .X(_05616_));
 sky130_fd_sc_hd__o311a_1 _13102_ (.A1(_05459_),
    .A2(_05461_),
    .A3(_05462_),
    .B1(_05614_),
    .C1(_05616_),
    .X(_05617_));
 sky130_fd_sc_hd__inv_2 _13103_ (.A(_04032_),
    .Y(_05618_));
 sky130_fd_sc_hd__o31a_2 _13104_ (.A1(_05609_),
    .A2(_05615_),
    .A3(_05617_),
    .B1(_05618_),
    .X(_05619_));
 sky130_fd_sc_hd__xnor2_4 _13105_ (.A(_04028_),
    .B(_05619_),
    .Y(_05620_));
 sky130_fd_sc_hd__and2_1 _13106_ (.A(_05608_),
    .B(_05620_),
    .X(_05622_));
 sky130_fd_sc_hd__inv_2 _13107_ (.A(_05622_),
    .Y(_05623_));
 sky130_fd_sc_hd__nor2_1 _13108_ (.A(_05605_),
    .B(_05623_),
    .Y(_05624_));
 sky130_fd_sc_hd__or2b_1 _13109_ (.A(_05217_),
    .B_N(_05216_),
    .X(_05625_));
 sky130_fd_sc_hd__o21a_2 _13110_ (.A1(_05154_),
    .A2(_05625_),
    .B1(_05218_),
    .X(_05626_));
 sky130_fd_sc_hd__nand2_1 _13111_ (.A(_05605_),
    .B(_05623_),
    .Y(_05627_));
 sky130_fd_sc_hd__o21a_1 _13112_ (.A1(_05624_),
    .A2(_05626_),
    .B1(_05627_),
    .X(_05628_));
 sky130_fd_sc_hd__xor2_1 _13113_ (.A(_04601_),
    .B(_04628_),
    .X(_05629_));
 sky130_fd_sc_hd__xnor2_2 _13114_ (.A(_05315_),
    .B(_05629_),
    .Y(_05630_));
 sky130_fd_sc_hd__xor2_2 _13115_ (.A(_05628_),
    .B(_05630_),
    .X(_05631_));
 sky130_fd_sc_hd__o31a_1 _13116_ (.A1(_03456_),
    .A2(_03496_),
    .A3(_03625_),
    .B1(_03671_),
    .X(_05633_));
 sky130_fd_sc_hd__xnor2_2 _13117_ (.A(_03669_),
    .B(_05633_),
    .Y(_05634_));
 sky130_fd_sc_hd__o31a_2 _13118_ (.A1(_05609_),
    .A2(_05615_),
    .A3(_05617_),
    .B1(_04031_),
    .X(_05635_));
 sky130_fd_sc_hd__xnor2_4 _13119_ (.A(_04029_),
    .B(_05635_),
    .Y(_05636_));
 sky130_fd_sc_hd__nor2_1 _13120_ (.A(_05634_),
    .B(_05636_),
    .Y(_05637_));
 sky130_fd_sc_hd__xor2_2 _13121_ (.A(_05608_),
    .B(_05620_),
    .X(_05638_));
 sky130_fd_sc_hd__nand2_1 _13122_ (.A(_05637_),
    .B(_05638_),
    .Y(_05639_));
 sky130_fd_sc_hd__or3_1 _13123_ (.A(_05215_),
    .B(_05171_),
    .C(_05212_),
    .X(_05640_));
 sky130_fd_sc_hd__nand2_2 _13124_ (.A(_05216_),
    .B(_05640_),
    .Y(_05641_));
 sky130_fd_sc_hd__nor2_1 _13125_ (.A(_05637_),
    .B(_05638_),
    .Y(_05642_));
 sky130_fd_sc_hd__a21o_2 _13126_ (.A1(_05639_),
    .A2(_05641_),
    .B1(_05642_),
    .X(_05644_));
 sky130_fd_sc_hd__xnor2_2 _13127_ (.A(_05605_),
    .B(_05623_),
    .Y(_05645_));
 sky130_fd_sc_hd__xnor2_4 _13128_ (.A(_05626_),
    .B(_05645_),
    .Y(_05646_));
 sky130_fd_sc_hd__xnor2_4 _13129_ (.A(_05644_),
    .B(_05646_),
    .Y(_05647_));
 sky130_fd_sc_hd__and2_4 _13130_ (.A(_05631_),
    .B(_05647_),
    .X(_05648_));
 sky130_fd_sc_hd__xnor2_2 _13131_ (.A(_03626_),
    .B(_03671_),
    .Y(_05649_));
 sky130_fd_sc_hd__or4_1 _13132_ (.A(_05609_),
    .B(_05615_),
    .C(_05617_),
    .D(_04031_),
    .X(_05650_));
 sky130_fd_sc_hd__or2b_4 _13133_ (.A(_05635_),
    .B_N(_05650_),
    .X(_05651_));
 sky130_fd_sc_hd__nor2_2 _13134_ (.A(_05649_),
    .B(_05651_),
    .Y(_05652_));
 sky130_fd_sc_hd__xor2_2 _13135_ (.A(_05634_),
    .B(_05636_),
    .X(_05653_));
 sky130_fd_sc_hd__nor2_1 _13136_ (.A(_05652_),
    .B(_05653_),
    .Y(_05655_));
 sky130_fd_sc_hd__o21a_1 _13137_ (.A1(_05182_),
    .A2(_05208_),
    .B1(_05211_),
    .X(_05656_));
 sky130_fd_sc_hd__a21oi_1 _13138_ (.A1(_05209_),
    .A2(_05210_),
    .B1(_05656_),
    .Y(_05657_));
 sky130_fd_sc_hd__nor2_1 _13139_ (.A(_05212_),
    .B(_05657_),
    .Y(_05658_));
 sky130_fd_sc_hd__a21oi_2 _13140_ (.A1(_05652_),
    .A2(_05653_),
    .B1(_05658_),
    .Y(_05659_));
 sky130_fd_sc_hd__nor2_2 _13141_ (.A(_05655_),
    .B(_05659_),
    .Y(_05660_));
 sky130_fd_sc_hd__xnor2_2 _13142_ (.A(_05637_),
    .B(_05638_),
    .Y(_05661_));
 sky130_fd_sc_hd__xnor2_4 _13143_ (.A(_05641_),
    .B(_05661_),
    .Y(_05662_));
 sky130_fd_sc_hd__xnor2_4 _13144_ (.A(_05660_),
    .B(_05662_),
    .Y(_05663_));
 sky130_fd_sc_hd__or2_1 _13145_ (.A(_05652_),
    .B(_05653_),
    .X(_05664_));
 sky130_fd_sc_hd__xnor2_1 _13146_ (.A(_05652_),
    .B(_05653_),
    .Y(_05666_));
 sky130_fd_sc_hd__a22o_1 _13147_ (.A1(_05664_),
    .A2(_05659_),
    .B1(_05666_),
    .B2(_05658_),
    .X(_05667_));
 sky130_fd_sc_hd__xor2_2 _13148_ (.A(_05649_),
    .B(_05651_),
    .X(_05668_));
 sky130_fd_sc_hd__xnor2_2 _13149_ (.A(_03053_),
    .B(_04624_),
    .Y(_05669_));
 sky130_fd_sc_hd__xnor2_4 _13150_ (.A(_04025_),
    .B(_04595_),
    .Y(_05670_));
 sky130_fd_sc_hd__and2_4 _13151_ (.A(_05669_),
    .B(_05670_),
    .X(_05671_));
 sky130_fd_sc_hd__inv_2 _13152_ (.A(_05182_),
    .Y(_05672_));
 sky130_fd_sc_hd__nand2_2 _13153_ (.A(_05211_),
    .B(_05672_),
    .Y(_05673_));
 sky130_fd_sc_hd__xnor2_4 _13154_ (.A(_05208_),
    .B(_05673_),
    .Y(_05674_));
 sky130_fd_sc_hd__a21o_1 _13155_ (.A1(_05668_),
    .A2(_05671_),
    .B1(_05674_),
    .X(_05675_));
 sky130_fd_sc_hd__o21a_1 _13156_ (.A1(_05668_),
    .A2(_05671_),
    .B1(_05675_),
    .X(_05677_));
 sky130_fd_sc_hd__xor2_2 _13157_ (.A(_05667_),
    .B(_05677_),
    .X(_05678_));
 sky130_fd_sc_hd__and2_4 _13158_ (.A(_05663_),
    .B(_05678_),
    .X(_05679_));
 sky130_fd_sc_hd__nand2_1 _13159_ (.A(_05648_),
    .B(_05679_),
    .Y(_05680_));
 sky130_fd_sc_hd__xnor2_2 _13160_ (.A(_05668_),
    .B(_05671_),
    .Y(_05681_));
 sky130_fd_sc_hd__xor2_4 _13161_ (.A(_05674_),
    .B(_05681_),
    .X(_05682_));
 sky130_fd_sc_hd__xnor2_2 _13162_ (.A(_05669_),
    .B(_05670_),
    .Y(_05683_));
 sky130_fd_sc_hd__a21oi_2 _13163_ (.A1(_05465_),
    .A2(_03624_),
    .B1(_03490_),
    .Y(_05684_));
 sky130_fd_sc_hd__xnor2_4 _13164_ (.A(_03493_),
    .B(_05684_),
    .Y(_05685_));
 sky130_fd_sc_hd__a21oi_2 _13165_ (.A1(_05616_),
    .A2(_05463_),
    .B1(_05612_),
    .Y(_05686_));
 sky130_fd_sc_hd__xnor2_4 _13166_ (.A(_04546_),
    .B(_05686_),
    .Y(_05688_));
 sky130_fd_sc_hd__or2_1 _13167_ (.A(_05685_),
    .B(_05688_),
    .X(_05689_));
 sky130_fd_sc_hd__or2_1 _13168_ (.A(_05683_),
    .B(_05689_),
    .X(_05690_));
 sky130_fd_sc_hd__xnor2_4 _13169_ (.A(_05196_),
    .B(_05206_),
    .Y(_05691_));
 sky130_fd_sc_hd__and2_1 _13170_ (.A(_05683_),
    .B(_05689_),
    .X(_05692_));
 sky130_fd_sc_hd__a21o_2 _13171_ (.A1(_05690_),
    .A2(_05691_),
    .B1(_05692_),
    .X(_05693_));
 sky130_fd_sc_hd__xor2_4 _13172_ (.A(_05682_),
    .B(_05693_),
    .X(_05694_));
 sky130_fd_sc_hd__xor2_2 _13173_ (.A(_05683_),
    .B(_05689_),
    .X(_05695_));
 sky130_fd_sc_hd__xnor2_4 _13174_ (.A(_05691_),
    .B(_05695_),
    .Y(_05696_));
 sky130_fd_sc_hd__nand3_1 _13175_ (.A(_03613_),
    .B(_03623_),
    .C(_04616_),
    .Y(_05697_));
 sky130_fd_sc_hd__o311a_1 _13176_ (.A1(_05479_),
    .A2(_04608_),
    .A3(_04611_),
    .B1(_05697_),
    .C1(_04621_),
    .X(_05699_));
 sky130_fd_sc_hd__xnor2_2 _13177_ (.A(_03622_),
    .B(_05699_),
    .Y(_05700_));
 sky130_fd_sc_hd__nand2_1 _13178_ (.A(_04403_),
    .B(_04454_),
    .Y(_05701_));
 sky130_fd_sc_hd__nand3_1 _13179_ (.A(_04531_),
    .B(_04536_),
    .C(_04490_),
    .Y(_05702_));
 sky130_fd_sc_hd__o311a_2 _13180_ (.A1(_05482_),
    .A2(_05701_),
    .A3(_04537_),
    .B1(_05702_),
    .C1(_04591_),
    .X(_05703_));
 sky130_fd_sc_hd__xnor2_4 _13181_ (.A(_04551_),
    .B(_05703_),
    .Y(_05704_));
 sky130_fd_sc_hd__and2_2 _13182_ (.A(_05700_),
    .B(_05704_),
    .X(_05705_));
 sky130_fd_sc_hd__xor2_4 _13183_ (.A(_05685_),
    .B(_05688_),
    .X(_05706_));
 sky130_fd_sc_hd__nand2_1 _13184_ (.A(_05202_),
    .B(_05205_),
    .Y(_05707_));
 sky130_fd_sc_hd__and2_1 _13185_ (.A(_05206_),
    .B(_05707_),
    .X(_05708_));
 sky130_fd_sc_hd__a21o_1 _13186_ (.A1(_05705_),
    .A2(_05706_),
    .B1(_05708_),
    .X(_05710_));
 sky130_fd_sc_hd__o21ai_4 _13187_ (.A1(_05705_),
    .A2(_05706_),
    .B1(_05710_),
    .Y(_05711_));
 sky130_fd_sc_hd__xnor2_4 _13188_ (.A(_05696_),
    .B(_05711_),
    .Y(_05712_));
 sky130_fd_sc_hd__nand2_1 _13189_ (.A(_05694_),
    .B(_05712_),
    .Y(_05713_));
 sky130_fd_sc_hd__xnor2_1 _13190_ (.A(_05705_),
    .B(_05706_),
    .Y(_05714_));
 sky130_fd_sc_hd__xnor2_2 _13191_ (.A(_05708_),
    .B(_05714_),
    .Y(_05715_));
 sky130_fd_sc_hd__nand2_1 _13192_ (.A(_05464_),
    .B(_05466_),
    .Y(_05716_));
 sky130_fd_sc_hd__inv_2 _13193_ (.A(_05716_),
    .Y(_05717_));
 sky130_fd_sc_hd__xor2_2 _13194_ (.A(_05700_),
    .B(_05704_),
    .X(_05718_));
 sky130_fd_sc_hd__nand2_1 _13195_ (.A(_05717_),
    .B(_05718_),
    .Y(_05719_));
 sky130_fd_sc_hd__nand2_1 _13196_ (.A(_05198_),
    .B(_05200_),
    .Y(_05721_));
 sky130_fd_sc_hd__xnor2_2 _13197_ (.A(_05199_),
    .B(_05721_),
    .Y(_05722_));
 sky130_fd_sc_hd__nor2_1 _13198_ (.A(_05717_),
    .B(_05718_),
    .Y(_05723_));
 sky130_fd_sc_hd__a21oi_2 _13199_ (.A1(_05719_),
    .A2(_05722_),
    .B1(_05723_),
    .Y(_05724_));
 sky130_fd_sc_hd__xor2_2 _13200_ (.A(_05715_),
    .B(_05724_),
    .X(_05725_));
 sky130_fd_sc_hd__and2_1 _13201_ (.A(_05457_),
    .B(_05469_),
    .X(_05726_));
 sky130_fd_sc_hd__or2_1 _13202_ (.A(_05457_),
    .B(_05469_),
    .X(_05727_));
 sky130_fd_sc_hd__o21ai_2 _13203_ (.A1(_05455_),
    .A2(_05726_),
    .B1(_05727_),
    .Y(_05728_));
 sky130_fd_sc_hd__xnor2_1 _13204_ (.A(_05717_),
    .B(_05718_),
    .Y(_05729_));
 sky130_fd_sc_hd__xnor2_2 _13205_ (.A(_05722_),
    .B(_05729_),
    .Y(_05730_));
 sky130_fd_sc_hd__xor2_2 _13206_ (.A(_05728_),
    .B(_05730_),
    .X(_05732_));
 sky130_fd_sc_hd__nand2_1 _13207_ (.A(_05725_),
    .B(_05732_),
    .Y(_05733_));
 sky130_fd_sc_hd__nand2_1 _13208_ (.A(_05715_),
    .B(_05724_),
    .Y(_05734_));
 sky130_fd_sc_hd__or2_1 _13209_ (.A(_05728_),
    .B(_05730_),
    .X(_05735_));
 sky130_fd_sc_hd__nor2_1 _13210_ (.A(_05715_),
    .B(_05724_),
    .Y(_05736_));
 sky130_fd_sc_hd__a21o_1 _13211_ (.A1(_05734_),
    .A2(_05735_),
    .B1(_05736_),
    .X(_05737_));
 sky130_fd_sc_hd__or2_1 _13212_ (.A(_05682_),
    .B(_05693_),
    .X(_05738_));
 sky130_fd_sc_hd__or2b_1 _13213_ (.A(_05711_),
    .B_N(_05696_),
    .X(_05739_));
 sky130_fd_sc_hd__and2_1 _13214_ (.A(_05682_),
    .B(_05693_),
    .X(_05740_));
 sky130_fd_sc_hd__a21oi_1 _13215_ (.A1(_05738_),
    .A2(_05739_),
    .B1(_05740_),
    .Y(_05741_));
 sky130_fd_sc_hd__o21ba_1 _13216_ (.A1(_05713_),
    .A2(_05737_),
    .B1_N(_05741_),
    .X(_05743_));
 sky130_fd_sc_hd__or3_1 _13217_ (.A(_05655_),
    .B(_05659_),
    .C(_05662_),
    .X(_05744_));
 sky130_fd_sc_hd__nand2_1 _13218_ (.A(_05667_),
    .B(_05677_),
    .Y(_05745_));
 sky130_fd_sc_hd__and2b_1 _13219_ (.A_N(_05660_),
    .B(_05662_),
    .X(_05746_));
 sky130_fd_sc_hd__a21oi_1 _13220_ (.A1(_05744_),
    .A2(_05745_),
    .B1(_05746_),
    .Y(_05747_));
 sky130_fd_sc_hd__inv_2 _13221_ (.A(_05644_),
    .Y(_05748_));
 sky130_fd_sc_hd__a22o_1 _13222_ (.A1(_05628_),
    .A2(_05630_),
    .B1(_05748_),
    .B2(_05646_),
    .X(_05749_));
 sky130_fd_sc_hd__o21a_1 _13223_ (.A1(_05628_),
    .A2(_05630_),
    .B1(_05749_),
    .X(_05750_));
 sky130_fd_sc_hd__a21o_1 _13224_ (.A1(_05648_),
    .A2(_05747_),
    .B1(_05750_),
    .X(_05751_));
 sky130_fd_sc_hd__o21ba_1 _13225_ (.A1(_05680_),
    .A2(_05743_),
    .B1_N(_05751_),
    .X(_05752_));
 sky130_fd_sc_hd__o41a_1 _13226_ (.A1(_05604_),
    .A2(_05680_),
    .A3(_05713_),
    .A4(_05733_),
    .B1(_05752_),
    .X(_05754_));
 sky130_fd_sc_hd__xor2_1 _13227_ (.A(_05424_),
    .B(_05754_),
    .X(net107));
 sky130_fd_sc_hd__o21ba_1 _13228_ (.A1(_05528_),
    .A2(_05582_),
    .B1_N(_05586_),
    .X(_05755_));
 sky130_fd_sc_hd__xnor2_4 _13229_ (.A(_05579_),
    .B(_05755_),
    .Y(net90));
 sky130_fd_sc_hd__and3_1 _13230_ (.A(_02713_),
    .B(_02714_),
    .C(_05579_),
    .X(_05756_));
 sky130_fd_sc_hd__o21a_1 _13231_ (.A1(_05590_),
    .A2(_02711_),
    .B1(_05578_),
    .X(_05757_));
 sky130_fd_sc_hd__a41o_1 _13232_ (.A1(_02716_),
    .A2(_02713_),
    .A3(_02715_),
    .A4(_05579_),
    .B1(_05757_),
    .X(_05758_));
 sky130_fd_sc_hd__a21oi_2 _13233_ (.A1(_02278_),
    .A2(_05756_),
    .B1(_05758_),
    .Y(_05759_));
 sky130_fd_sc_hd__xnor2_4 _13234_ (.A(_05575_),
    .B(_05759_),
    .Y(net91));
 sky130_fd_sc_hd__a32o_1 _13235_ (.A1(_05575_),
    .A2(_05579_),
    .A3(_05585_),
    .B1(_05591_),
    .B2(_05589_),
    .X(_05760_));
 sky130_fd_sc_hd__inv_2 _13236_ (.A(_05760_),
    .Y(_05762_));
 sky130_fd_sc_hd__and4_1 _13237_ (.A(_02491_),
    .B(_02713_),
    .C(_05575_),
    .D(_05579_),
    .X(_05763_));
 sky130_fd_sc_hd__nand2_1 _13238_ (.A(_02494_),
    .B(_05763_),
    .Y(_05764_));
 sky130_fd_sc_hd__nand4_2 _13239_ (.A(_01640_),
    .B(_02046_),
    .C(_02492_),
    .D(_05763_),
    .Y(_05765_));
 sky130_fd_sc_hd__and3_1 _13240_ (.A(_05762_),
    .B(_05764_),
    .C(_05765_),
    .X(_05766_));
 sky130_fd_sc_hd__xnor2_4 _13241_ (.A(_05562_),
    .B(_05766_),
    .Y(net92));
 sky130_fd_sc_hd__nand3_1 _13242_ (.A(_05572_),
    .B(_05568_),
    .C(_05570_),
    .Y(_05767_));
 sky130_fd_sc_hd__and3b_2 _13243_ (.A_N(_05573_),
    .B(_05767_),
    .C(_05562_),
    .X(_05768_));
 sky130_fd_sc_hd__and3_1 _13244_ (.A(_02713_),
    .B(_05579_),
    .C(_05768_),
    .X(_05769_));
 sky130_fd_sc_hd__and3_1 _13245_ (.A(_05548_),
    .B(_05557_),
    .C(_05560_),
    .X(_05770_));
 sky130_fd_sc_hd__a21oi_2 _13246_ (.A1(_05592_),
    .A2(_05767_),
    .B1(_05770_),
    .Y(_05772_));
 sky130_fd_sc_hd__a221oi_4 _13247_ (.A1(_05757_),
    .A2(_05768_),
    .B1(_05769_),
    .B2(_02717_),
    .C1(_05772_),
    .Y(_05773_));
 sky130_fd_sc_hd__nand4_1 _13248_ (.A(_01837_),
    .B(_02045_),
    .C(_02274_),
    .D(_02491_),
    .Y(_05774_));
 sky130_fd_sc_hd__nand3_1 _13249_ (.A(_02713_),
    .B(_05579_),
    .C(_05768_),
    .Y(_05775_));
 sky130_fd_sc_hd__a211o_4 _13250_ (.A1(_01647_),
    .A2(_01648_),
    .B1(_05774_),
    .C1(_05775_),
    .X(_05776_));
 sky130_fd_sc_hd__and2_4 _13251_ (.A(_05776_),
    .B(_05773_),
    .X(_05777_));
 sky130_fd_sc_hd__xnor2_2 _13252_ (.A(_05546_),
    .B(_05777_),
    .Y(net93));
 sky130_fd_sc_hd__xor2_4 _13253_ (.A(_05524_),
    .B(net130),
    .X(net94));
 sky130_fd_sc_hd__or2b_2 _13254_ (.A(_05505_),
    .B_N(_05506_),
    .X(_05778_));
 sky130_fd_sc_hd__and2_1 _13255_ (.A(_05524_),
    .B(_05546_),
    .X(_05779_));
 sky130_fd_sc_hd__and2_1 _13256_ (.A(_05768_),
    .B(_05779_),
    .X(_05781_));
 sky130_fd_sc_hd__and2_1 _13257_ (.A(_05758_),
    .B(_05781_),
    .X(_05782_));
 sky130_fd_sc_hd__and2_1 _13258_ (.A(_05519_),
    .B(_05523_),
    .X(_05783_));
 sky130_fd_sc_hd__a21oi_2 _13259_ (.A1(_05596_),
    .A2(_05545_),
    .B1(_05783_),
    .Y(_05784_));
 sky130_fd_sc_hd__a21o_1 _13260_ (.A1(_05772_),
    .A2(_05779_),
    .B1(_05784_),
    .X(_05785_));
 sky130_fd_sc_hd__a311o_4 _13261_ (.A1(_02278_),
    .A2(_05756_),
    .A3(_05781_),
    .B1(_05782_),
    .C1(_05785_),
    .X(_05786_));
 sky130_fd_sc_hd__xnor2_4 _13262_ (.A(_05778_),
    .B(_05786_),
    .Y(net95));
 sky130_fd_sc_hd__xnor2_4 _13263_ (.A(_05474_),
    .B(_05490_),
    .Y(_05787_));
 sky130_fd_sc_hd__and3_1 _13264_ (.A(_05507_),
    .B(_05524_),
    .C(_05563_),
    .X(_05788_));
 sky130_fd_sc_hd__a31o_1 _13265_ (.A1(_05507_),
    .A2(_05524_),
    .A3(_05593_),
    .B1(_05597_),
    .X(_05789_));
 sky130_fd_sc_hd__a21o_1 _13266_ (.A1(_05760_),
    .A2(_05788_),
    .B1(_05789_),
    .X(_05791_));
 sky130_fd_sc_hd__a31o_4 _13267_ (.A1(_02495_),
    .A2(_05763_),
    .A3(_05788_),
    .B1(_05791_),
    .X(_05792_));
 sky130_fd_sc_hd__xnor2_4 _13268_ (.A(_05787_),
    .B(_05792_),
    .Y(net96));
 sky130_fd_sc_hd__nor2_1 _13269_ (.A(_05787_),
    .B(_05778_),
    .Y(_05793_));
 sky130_fd_sc_hd__nand2_1 _13270_ (.A(_05779_),
    .B(_05793_),
    .Y(_05794_));
 sky130_fd_sc_hd__a21o_1 _13271_ (.A1(_05773_),
    .A2(_05776_),
    .B1(_05794_),
    .X(_05795_));
 sky130_fd_sc_hd__and2_1 _13272_ (.A(_05474_),
    .B(_05490_),
    .X(_05796_));
 sky130_fd_sc_hd__a21oi_1 _13273_ (.A1(_05600_),
    .A2(_05506_),
    .B1(_05796_),
    .Y(_05797_));
 sky130_fd_sc_hd__a21oi_2 _13274_ (.A1(_05784_),
    .A2(_05793_),
    .B1(_05797_),
    .Y(_05798_));
 sky130_fd_sc_hd__nand2_2 _13275_ (.A(_05795_),
    .B(_05798_),
    .Y(_05799_));
 sky130_fd_sc_hd__xor2_4 _13276_ (.A(_05472_),
    .B(_05799_),
    .X(net97));
 sky130_fd_sc_hd__xnor2_1 _13277_ (.A(_05604_),
    .B(_05732_),
    .Y(net99));
 sky130_fd_sc_hd__and2_1 _13278_ (.A(_05472_),
    .B(_05732_),
    .X(_05801_));
 sky130_fd_sc_hd__and2_1 _13279_ (.A(_05793_),
    .B(_05801_),
    .X(_05802_));
 sky130_fd_sc_hd__and2_1 _13280_ (.A(_05728_),
    .B(_05730_),
    .X(_05803_));
 sky130_fd_sc_hd__a21oi_1 _13281_ (.A1(_05598_),
    .A2(_05735_),
    .B1(_05803_),
    .Y(_05804_));
 sky130_fd_sc_hd__a21o_1 _13282_ (.A1(_05797_),
    .A2(_05801_),
    .B1(_05804_),
    .X(_05805_));
 sky130_fd_sc_hd__a21oi_1 _13283_ (.A1(_05786_),
    .A2(_05802_),
    .B1(_05805_),
    .Y(_05806_));
 sky130_fd_sc_hd__xnor2_1 _13284_ (.A(_05725_),
    .B(_05806_),
    .Y(net100));
 sky130_fd_sc_hd__and4_2 _13285_ (.A(_05472_),
    .B(_05491_),
    .C(_05725_),
    .D(_05732_),
    .X(_05807_));
 sky130_fd_sc_hd__nand2_1 _13286_ (.A(_05788_),
    .B(_05807_),
    .Y(_05809_));
 sky130_fd_sc_hd__a31o_2 _13287_ (.A1(_05762_),
    .A2(_05764_),
    .A3(_05765_),
    .B1(_05809_),
    .X(_05810_));
 sky130_fd_sc_hd__o21a_1 _13288_ (.A1(_05602_),
    .A2(_05733_),
    .B1(_05737_),
    .X(_05811_));
 sky130_fd_sc_hd__nand2_1 _13289_ (.A(_05789_),
    .B(_05807_),
    .Y(_05812_));
 sky130_fd_sc_hd__nand3_2 _13290_ (.A(_05810_),
    .B(_05811_),
    .C(_05812_),
    .Y(_05813_));
 sky130_fd_sc_hd__xor2_4 _13291_ (.A(_05712_),
    .B(_05813_),
    .X(net101));
 sky130_fd_sc_hd__and2_1 _13292_ (.A(_05712_),
    .B(_05725_),
    .X(_05814_));
 sky130_fd_sc_hd__nand2_1 _13293_ (.A(_05801_),
    .B(_05814_),
    .Y(_05815_));
 sky130_fd_sc_hd__or2_1 _13294_ (.A(_05798_),
    .B(_05815_),
    .X(_05816_));
 sky130_fd_sc_hd__and2b_1 _13295_ (.A_N(_05696_),
    .B(_05711_),
    .X(_05817_));
 sky130_fd_sc_hd__a21oi_2 _13296_ (.A1(_05739_),
    .A2(_05734_),
    .B1(_05817_),
    .Y(_05819_));
 sky130_fd_sc_hd__a21oi_2 _13297_ (.A1(_05804_),
    .A2(_05814_),
    .B1(_05819_),
    .Y(_05820_));
 sky130_fd_sc_hd__o311a_4 _13298_ (.A1(_05777_),
    .A2(_05794_),
    .A3(_05815_),
    .B1(_05816_),
    .C1(_05820_),
    .X(_05821_));
 sky130_fd_sc_hd__xnor2_4 _13299_ (.A(_05694_),
    .B(_05821_),
    .Y(net102));
 sky130_fd_sc_hd__nor2_1 _13300_ (.A(_05713_),
    .B(_05733_),
    .Y(_05822_));
 sky130_fd_sc_hd__inv_2 _13301_ (.A(_05743_),
    .Y(_05823_));
 sky130_fd_sc_hd__and2_1 _13302_ (.A(_05603_),
    .B(_05822_),
    .X(_05824_));
 sky130_fd_sc_hd__a311o_4 _13303_ (.A1(_05525_),
    .A2(_05595_),
    .A3(_05822_),
    .B1(_05823_),
    .C1(_05824_),
    .X(_05825_));
 sky130_fd_sc_hd__xor2_2 _13304_ (.A(_05678_),
    .B(_05825_),
    .X(net103));
 sky130_fd_sc_hd__and2_1 _13305_ (.A(_05678_),
    .B(_05694_),
    .X(_05826_));
 sky130_fd_sc_hd__nor2_1 _13306_ (.A(_05667_),
    .B(_05677_),
    .Y(_05828_));
 sky130_fd_sc_hd__a21oi_1 _13307_ (.A1(_05745_),
    .A2(_05738_),
    .B1(_05828_),
    .Y(_05829_));
 sky130_fd_sc_hd__a21o_1 _13308_ (.A1(_05819_),
    .A2(_05826_),
    .B1(_05829_),
    .X(_05830_));
 sky130_fd_sc_hd__and2_1 _13309_ (.A(_05814_),
    .B(_05826_),
    .X(_05831_));
 sky130_fd_sc_hd__and2_1 _13310_ (.A(_05805_),
    .B(_05831_),
    .X(_05832_));
 sky130_fd_sc_hd__a31o_2 _13311_ (.A1(_05786_),
    .A2(_05802_),
    .A3(_05831_),
    .B1(_05832_),
    .X(_05833_));
 sky130_fd_sc_hd__nor2_1 _13312_ (.A(_05830_),
    .B(_05833_),
    .Y(_05834_));
 sky130_fd_sc_hd__xnor2_2 _13313_ (.A(_05663_),
    .B(_05834_),
    .Y(net104));
 sky130_fd_sc_hd__nand3_1 _13314_ (.A(_05679_),
    .B(_05694_),
    .C(_05712_),
    .Y(_05835_));
 sky130_fd_sc_hd__inv_2 _13315_ (.A(_05835_),
    .Y(_05836_));
 sky130_fd_sc_hd__nor2_1 _13316_ (.A(_05811_),
    .B(_05835_),
    .Y(_05838_));
 sky130_fd_sc_hd__a21oi_1 _13317_ (.A1(_05679_),
    .A2(_05741_),
    .B1(_05747_),
    .Y(_05839_));
 sky130_fd_sc_hd__inv_2 _13318_ (.A(_05839_),
    .Y(_05840_));
 sky130_fd_sc_hd__a311o_4 _13319_ (.A1(_05792_),
    .A2(_05807_),
    .A3(_05836_),
    .B1(_05838_),
    .C1(_05840_),
    .X(_05841_));
 sky130_fd_sc_hd__xor2_4 _13320_ (.A(_05647_),
    .B(_05841_),
    .X(net105));
 sky130_fd_sc_hd__nand3_2 _13321_ (.A(_05647_),
    .B(_05663_),
    .C(_05826_),
    .Y(_05842_));
 sky130_fd_sc_hd__a211o_1 _13322_ (.A1(_05795_),
    .A2(_05798_),
    .B1(_05815_),
    .C1(_05842_),
    .X(_05843_));
 sky130_fd_sc_hd__nand2_1 _13323_ (.A(_05748_),
    .B(_05646_),
    .Y(_05844_));
 sky130_fd_sc_hd__nor2_1 _13324_ (.A(_05748_),
    .B(_05646_),
    .Y(_05845_));
 sky130_fd_sc_hd__a21oi_1 _13325_ (.A1(_05844_),
    .A2(_05744_),
    .B1(_05845_),
    .Y(_05846_));
 sky130_fd_sc_hd__a31o_1 _13326_ (.A1(_05647_),
    .A2(_05663_),
    .A3(_05829_),
    .B1(_05846_),
    .X(_05848_));
 sky130_fd_sc_hd__o21ba_1 _13327_ (.A1(_05820_),
    .A2(_05842_),
    .B1_N(_05848_),
    .X(_05849_));
 sky130_fd_sc_hd__nand2_1 _13328_ (.A(_05843_),
    .B(_05849_),
    .Y(_05850_));
 sky130_fd_sc_hd__xor2_1 _13329_ (.A(_05631_),
    .B(_05850_),
    .X(net106));
 sky130_fd_sc_hd__and2b_1 _13330_ (.A_N(_05318_),
    .B(_05419_),
    .X(_05851_));
 sky130_fd_sc_hd__or2b_1 _13331_ (.A(_05411_),
    .B_N(_05415_),
    .X(_05852_));
 sky130_fd_sc_hd__and2b_1 _13332_ (.A_N(_05362_),
    .B(_05408_),
    .X(_05853_));
 sky130_fd_sc_hd__nand2_1 _13333_ (.A(_05325_),
    .B(_05332_),
    .Y(_05854_));
 sky130_fd_sc_hd__o21ba_1 _13334_ (.A1(_05327_),
    .A2(_05330_),
    .B1_N(_05328_),
    .X(_05855_));
 sky130_fd_sc_hd__a22o_1 _13335_ (.A1(_00745_),
    .A2(_02724_),
    .B1(_02728_),
    .B2(_00914_),
    .X(_05856_));
 sky130_fd_sc_hd__nand4_1 _13336_ (.A(_00914_),
    .B(_00745_),
    .C(_02724_),
    .D(_02728_),
    .Y(_05858_));
 sky130_fd_sc_hd__nand2_1 _13337_ (.A(_05856_),
    .B(_05858_),
    .Y(_05859_));
 sky130_fd_sc_hd__xor2_1 _13338_ (.A(_05855_),
    .B(_05859_),
    .X(_05860_));
 sky130_fd_sc_hd__and3_1 _13339_ (.A(_05326_),
    .B(_05331_),
    .C(_05860_),
    .X(_05861_));
 sky130_fd_sc_hd__and2_1 _13340_ (.A(_05326_),
    .B(_05331_),
    .X(_05862_));
 sky130_fd_sc_hd__nor2_1 _13341_ (.A(_05862_),
    .B(_05860_),
    .Y(_05863_));
 sky130_fd_sc_hd__or2_1 _13342_ (.A(_05861_),
    .B(_05863_),
    .X(_05864_));
 sky130_fd_sc_hd__and3_1 _13343_ (.A(_05854_),
    .B(_05336_),
    .C(_05864_),
    .X(_05865_));
 sky130_fd_sc_hd__a21oi_1 _13344_ (.A1(_05854_),
    .A2(_05336_),
    .B1(_05864_),
    .Y(_05866_));
 sky130_fd_sc_hd__nor2_1 _13345_ (.A(_05865_),
    .B(_05866_),
    .Y(_05867_));
 sky130_fd_sc_hd__nand2_1 _13346_ (.A(_05340_),
    .B(_05348_),
    .Y(_05869_));
 sky130_fd_sc_hd__o21ba_1 _13347_ (.A1(_05342_),
    .A2(_05345_),
    .B1_N(_05343_),
    .X(_05870_));
 sky130_fd_sc_hd__a22o_1 _13348_ (.A1(_01584_),
    .A2(_02306_),
    .B1(_02305_),
    .B2(_01586_),
    .X(_05871_));
 sky130_fd_sc_hd__nand4_1 _13349_ (.A(_01600_),
    .B(_01585_),
    .C(_02306_),
    .D(_02857_),
    .Y(_05872_));
 sky130_fd_sc_hd__nand2_1 _13350_ (.A(_05871_),
    .B(_05872_),
    .Y(_05873_));
 sky130_fd_sc_hd__xor2_1 _13351_ (.A(_05870_),
    .B(_05873_),
    .X(_05874_));
 sky130_fd_sc_hd__and3_1 _13352_ (.A(_05341_),
    .B(_05347_),
    .C(_05874_),
    .X(_05875_));
 sky130_fd_sc_hd__and2_1 _13353_ (.A(_05341_),
    .B(_05347_),
    .X(_05876_));
 sky130_fd_sc_hd__nor2_1 _13354_ (.A(_05876_),
    .B(_05874_),
    .Y(_05877_));
 sky130_fd_sc_hd__or2_1 _13355_ (.A(_05875_),
    .B(_05877_),
    .X(_05878_));
 sky130_fd_sc_hd__and3_1 _13356_ (.A(_05869_),
    .B(_05351_),
    .C(_05878_),
    .X(_05880_));
 sky130_fd_sc_hd__a21oi_1 _13357_ (.A1(_05869_),
    .A2(_05351_),
    .B1(_05878_),
    .Y(_05881_));
 sky130_fd_sc_hd__nor2_1 _13358_ (.A(_05880_),
    .B(_05881_),
    .Y(_05882_));
 sky130_fd_sc_hd__xor2_1 _13359_ (.A(_05867_),
    .B(_05882_),
    .X(_05883_));
 sky130_fd_sc_hd__a21oi_1 _13360_ (.A1(_05337_),
    .A2(_05352_),
    .B1(_05883_),
    .Y(_05884_));
 sky130_fd_sc_hd__nand3_1 _13361_ (.A(_05337_),
    .B(_05352_),
    .C(_05883_),
    .Y(_05885_));
 sky130_fd_sc_hd__or2b_1 _13362_ (.A(_05884_),
    .B_N(_05885_),
    .X(_05886_));
 sky130_fd_sc_hd__and3_1 _13363_ (.A(_00416_),
    .B(_01288_),
    .C(_02720_),
    .X(_05887_));
 sky130_fd_sc_hd__a22o_1 _13364_ (.A1(_01289_),
    .A2(_02759_),
    .B1(_02721_),
    .B2(_02008_),
    .X(_05888_));
 sky130_fd_sc_hd__a21bo_1 _13365_ (.A1(_02765_),
    .A2(_05887_),
    .B1_N(_05888_),
    .X(_05889_));
 sky130_fd_sc_hd__xnor2_1 _13366_ (.A(_05886_),
    .B(_05889_),
    .Y(_05891_));
 sky130_fd_sc_hd__a21o_1 _13367_ (.A1(_05292_),
    .A2(_05354_),
    .B1(_05353_),
    .X(_05892_));
 sky130_fd_sc_hd__a32o_1 _13368_ (.A1(_05292_),
    .A2(_05353_),
    .A3(_05354_),
    .B1(_02765_),
    .B2(_02008_),
    .X(_05893_));
 sky130_fd_sc_hd__nand2_1 _13369_ (.A(_05892_),
    .B(_05893_),
    .Y(_05894_));
 sky130_fd_sc_hd__xnor2_1 _13370_ (.A(_05891_),
    .B(_05894_),
    .Y(_05895_));
 sky130_fd_sc_hd__nand2_1 _13371_ (.A(_05360_),
    .B(_05895_),
    .Y(_05896_));
 sky130_fd_sc_hd__a211o_1 _13372_ (.A1(_05320_),
    .A2(_05321_),
    .B1(_05359_),
    .C1(_05895_),
    .X(_05897_));
 sky130_fd_sc_hd__and2_1 _13373_ (.A(_05896_),
    .B(_05897_),
    .X(_05898_));
 sky130_fd_sc_hd__nand2_1 _13374_ (.A(_05366_),
    .B(_05375_),
    .Y(_05899_));
 sky130_fd_sc_hd__and2_1 _13375_ (.A(_05367_),
    .B(_05374_),
    .X(_05900_));
 sky130_fd_sc_hd__a31oi_2 _13376_ (.A1(_00607_),
    .A2(_03744_),
    .A3(_05372_),
    .B1(_05371_),
    .Y(_05902_));
 sky130_fd_sc_hd__a22o_1 _13377_ (.A1(_01504_),
    .A2(_03738_),
    .B1(_03744_),
    .B2(_01508_),
    .X(_05903_));
 sky130_fd_sc_hd__nand4_1 _13378_ (.A(_01664_),
    .B(_01505_),
    .C(_03738_),
    .D(_03744_),
    .Y(_05904_));
 sky130_fd_sc_hd__nand2_1 _13379_ (.A(_05903_),
    .B(_05904_),
    .Y(_05905_));
 sky130_fd_sc_hd__xor2_1 _13380_ (.A(_05902_),
    .B(_05905_),
    .X(_05906_));
 sky130_fd_sc_hd__and2_1 _13381_ (.A(_05900_),
    .B(_05906_),
    .X(_05907_));
 sky130_fd_sc_hd__nor2_1 _13382_ (.A(_05900_),
    .B(_05906_),
    .Y(_05908_));
 sky130_fd_sc_hd__or2_1 _13383_ (.A(_05907_),
    .B(_05908_),
    .X(_05909_));
 sky130_fd_sc_hd__and3_1 _13384_ (.A(_05899_),
    .B(_05378_),
    .C(_05909_),
    .X(_05910_));
 sky130_fd_sc_hd__a21oi_1 _13385_ (.A1(_05899_),
    .A2(_05378_),
    .B1(_05909_),
    .Y(_05911_));
 sky130_fd_sc_hd__nor2_1 _13386_ (.A(_05910_),
    .B(_05911_),
    .Y(_05913_));
 sky130_fd_sc_hd__nand2_1 _13387_ (.A(_05383_),
    .B(_05392_),
    .Y(_05914_));
 sky130_fd_sc_hd__and2_1 _13388_ (.A(_05384_),
    .B(_05391_),
    .X(_05915_));
 sky130_fd_sc_hd__a31oi_2 _13389_ (.A1(_00375_),
    .A2(_02673_),
    .A3(_05388_),
    .B1(_05387_),
    .Y(_05916_));
 sky130_fd_sc_hd__a22o_1 _13390_ (.A1(_00779_),
    .A2(_03681_),
    .B1(_02673_),
    .B2(_01518_),
    .X(_05917_));
 sky130_fd_sc_hd__nand4_1 _13391_ (.A(_01518_),
    .B(_01517_),
    .C(_03681_),
    .D(_02673_),
    .Y(_05918_));
 sky130_fd_sc_hd__nand2_1 _13392_ (.A(_05917_),
    .B(_05918_),
    .Y(_05919_));
 sky130_fd_sc_hd__xor2_1 _13393_ (.A(_05916_),
    .B(_05919_),
    .X(_05920_));
 sky130_fd_sc_hd__and2_1 _13394_ (.A(_05915_),
    .B(_05920_),
    .X(_05921_));
 sky130_fd_sc_hd__nor2_1 _13395_ (.A(_05915_),
    .B(_05920_),
    .Y(_05922_));
 sky130_fd_sc_hd__or2_1 _13396_ (.A(_05921_),
    .B(_05922_),
    .X(_05924_));
 sky130_fd_sc_hd__and3_1 _13397_ (.A(_05914_),
    .B(_05395_),
    .C(_05924_),
    .X(_05925_));
 sky130_fd_sc_hd__a21oi_1 _13398_ (.A1(_05914_),
    .A2(_05395_),
    .B1(_05924_),
    .Y(_05926_));
 sky130_fd_sc_hd__nor2_1 _13399_ (.A(_05925_),
    .B(_05926_),
    .Y(_05927_));
 sky130_fd_sc_hd__xnor2_1 _13400_ (.A(_05913_),
    .B(_05927_),
    .Y(_05928_));
 sky130_fd_sc_hd__nand2_1 _13401_ (.A(_05397_),
    .B(_05928_),
    .Y(_05929_));
 sky130_fd_sc_hd__or2_1 _13402_ (.A(_05397_),
    .B(_05928_),
    .X(_05930_));
 sky130_fd_sc_hd__nand2_1 _13403_ (.A(_05929_),
    .B(_05930_),
    .Y(_05931_));
 sky130_fd_sc_hd__a22o_1 _13404_ (.A1(_03414_),
    .A2(_01956_),
    .B1(_03687_),
    .B2(_04714_),
    .X(_05932_));
 sky130_fd_sc_hd__and4_1 _13405_ (.A(_01066_),
    .B(_03414_),
    .C(_01955_),
    .D(_03686_),
    .X(_05933_));
 sky130_fd_sc_hd__inv_2 _13406_ (.A(_05933_),
    .Y(_05935_));
 sky130_fd_sc_hd__and2_1 _13407_ (.A(_05932_),
    .B(_05935_),
    .X(_05936_));
 sky130_fd_sc_hd__xor2_2 _13408_ (.A(_05931_),
    .B(_05936_),
    .X(_05937_));
 sky130_fd_sc_hd__a21o_1 _13409_ (.A1(_05248_),
    .A2(_05400_),
    .B1(_05399_),
    .X(_05938_));
 sky130_fd_sc_hd__a32o_1 _13410_ (.A1(_05248_),
    .A2(_05399_),
    .A3(_05400_),
    .B1(_01956_),
    .B2(_04714_),
    .X(_05939_));
 sky130_fd_sc_hd__nand2_1 _13411_ (.A(_05938_),
    .B(_05939_),
    .Y(_05940_));
 sky130_fd_sc_hd__xnor2_2 _13412_ (.A(_05937_),
    .B(_05940_),
    .Y(_05941_));
 sky130_fd_sc_hd__xnor2_2 _13413_ (.A(_05406_),
    .B(_05941_),
    .Y(_05942_));
 sky130_fd_sc_hd__nand2_1 _13414_ (.A(_05898_),
    .B(_05942_),
    .Y(_05943_));
 sky130_fd_sc_hd__or2_1 _13415_ (.A(_05898_),
    .B(_05942_),
    .X(_05944_));
 sky130_fd_sc_hd__and3_1 _13416_ (.A(_05853_),
    .B(_05943_),
    .C(_05944_),
    .X(_05946_));
 sky130_fd_sc_hd__a21oi_1 _13417_ (.A1(_05943_),
    .A2(_05944_),
    .B1(_05853_),
    .Y(_05947_));
 sky130_fd_sc_hd__or2_1 _13418_ (.A(_05946_),
    .B(_05947_),
    .X(_05948_));
 sky130_fd_sc_hd__a22o_1 _13419_ (.A1(_01183_),
    .A2(_01415_),
    .B1(_01252_),
    .B2(_01108_),
    .X(_05949_));
 sky130_fd_sc_hd__and4_1 _13420_ (.A(_01061_),
    .B(_01181_),
    .C(_01414_),
    .D(_01250_),
    .X(_05950_));
 sky130_fd_sc_hd__inv_2 _13421_ (.A(_05950_),
    .Y(_05951_));
 sky130_fd_sc_hd__and2_1 _13422_ (.A(_05949_),
    .B(_05951_),
    .X(_05952_));
 sky130_fd_sc_hd__xnor2_1 _13423_ (.A(_05948_),
    .B(_05952_),
    .Y(_05953_));
 sky130_fd_sc_hd__and3_1 _13424_ (.A(_05413_),
    .B(_05852_),
    .C(_05953_),
    .X(_05954_));
 sky130_fd_sc_hd__a21o_1 _13425_ (.A1(_05413_),
    .A2(_05852_),
    .B1(_05953_),
    .X(_05955_));
 sky130_fd_sc_hd__and2b_1 _13426_ (.A_N(_05954_),
    .B(_05955_),
    .X(_05957_));
 sky130_fd_sc_hd__xor2_2 _13427_ (.A(_05417_),
    .B(_05957_),
    .X(_05958_));
 sky130_fd_sc_hd__nand2_1 _13428_ (.A(_05851_),
    .B(_05957_),
    .Y(_05959_));
 sky130_fd_sc_hd__o21ai_4 _13429_ (.A1(_05851_),
    .A2(_05958_),
    .B1(_05959_),
    .Y(_05960_));
 sky130_fd_sc_hd__and2b_1 _13430_ (.A_N(_05424_),
    .B(_05631_),
    .X(_05961_));
 sky130_fd_sc_hd__and3_2 _13431_ (.A(_05647_),
    .B(_05663_),
    .C(_05961_),
    .X(_05962_));
 sky130_fd_sc_hd__a21o_1 _13432_ (.A1(_05628_),
    .A2(_05630_),
    .B1(_05421_),
    .X(_05963_));
 sky130_fd_sc_hd__and2_1 _13433_ (.A(_05422_),
    .B(_05963_),
    .X(_05964_));
 sky130_fd_sc_hd__a21o_1 _13434_ (.A1(_05846_),
    .A2(_05961_),
    .B1(_05964_),
    .X(_05965_));
 sky130_fd_sc_hd__a21o_1 _13435_ (.A1(_05830_),
    .A2(_05962_),
    .B1(_05965_),
    .X(_05966_));
 sky130_fd_sc_hd__a21oi_4 _13436_ (.A1(_05833_),
    .A2(_05962_),
    .B1(_05966_),
    .Y(_05968_));
 sky130_fd_sc_hd__xor2_4 _13437_ (.A(_05960_),
    .B(_05968_),
    .X(net108));
 sky130_fd_sc_hd__buf_2 _13438_ (.A(_03785_),
    .X(_05969_));
 sky130_fd_sc_hd__and4_1 _13439_ (.A(_01181_),
    .B(_01250_),
    .C(_02721_),
    .D(_02726_),
    .X(_05970_));
 sky130_fd_sc_hd__inv_2 _13440_ (.A(_05970_),
    .Y(_05971_));
 sky130_fd_sc_hd__a22o_1 _13441_ (.A1(_01250_),
    .A2(_02721_),
    .B1(_02735_),
    .B2(_01182_),
    .X(_05972_));
 sky130_fd_sc_hd__and4_1 _13442_ (.A(_05969_),
    .B(_02765_),
    .C(_05971_),
    .D(_05972_),
    .X(_05973_));
 sky130_fd_sc_hd__a22oi_1 _13443_ (.A1(_05969_),
    .A2(_02766_),
    .B1(_05971_),
    .B2(_05972_),
    .Y(_05974_));
 sky130_fd_sc_hd__nor2_1 _13444_ (.A(_05973_),
    .B(_05974_),
    .Y(_05975_));
 sky130_fd_sc_hd__and4_1 _13445_ (.A(_01183_),
    .B(_01252_),
    .C(_02766_),
    .D(_02722_),
    .X(_05976_));
 sky130_fd_sc_hd__nand2_1 _13446_ (.A(_05975_),
    .B(_05976_),
    .Y(_05978_));
 sky130_fd_sc_hd__and4_1 _13447_ (.A(_01182_),
    .B(_01252_),
    .C(_02735_),
    .D(_02731_),
    .X(_05979_));
 sky130_fd_sc_hd__a22o_1 _13448_ (.A1(_01252_),
    .A2(_02736_),
    .B1(_02731_),
    .B2(_01182_),
    .X(_05980_));
 sky130_fd_sc_hd__and2b_1 _13449_ (.A_N(_05979_),
    .B(_05980_),
    .X(_05981_));
 sky130_fd_sc_hd__nand2_1 _13450_ (.A(_05969_),
    .B(_02722_),
    .Y(_05982_));
 sky130_fd_sc_hd__xnor2_1 _13451_ (.A(_05981_),
    .B(_05982_),
    .Y(_05983_));
 sky130_fd_sc_hd__or2_1 _13452_ (.A(_05970_),
    .B(_05973_),
    .X(_05984_));
 sky130_fd_sc_hd__buf_2 _13453_ (.A(_03783_),
    .X(_05985_));
 sky130_fd_sc_hd__nand2_1 _13454_ (.A(_05985_),
    .B(_02766_),
    .Y(_05986_));
 sky130_fd_sc_hd__xnor2_1 _13455_ (.A(_05984_),
    .B(_05986_),
    .Y(_05987_));
 sky130_fd_sc_hd__nand2_1 _13456_ (.A(_05983_),
    .B(_05987_),
    .Y(_05989_));
 sky130_fd_sc_hd__or2_1 _13457_ (.A(_05983_),
    .B(_05987_),
    .X(_05990_));
 sky130_fd_sc_hd__nand2_1 _13458_ (.A(_05989_),
    .B(_05990_),
    .Y(_05991_));
 sky130_fd_sc_hd__nor2_1 _13459_ (.A(_05978_),
    .B(_05991_),
    .Y(_05992_));
 sky130_fd_sc_hd__or2b_1 _13460_ (.A(_05986_),
    .B_N(_05984_),
    .X(_05993_));
 sky130_fd_sc_hd__a31o_1 _13461_ (.A1(_05969_),
    .A2(_02722_),
    .A3(_05980_),
    .B1(_05979_),
    .X(_05994_));
 sky130_fd_sc_hd__nand2_1 _13462_ (.A(_05969_),
    .B(_02735_),
    .Y(_05995_));
 sky130_fd_sc_hd__a21boi_1 _13463_ (.A1(_01252_),
    .A2(_02737_),
    .B1_N(_05995_),
    .Y(_05996_));
 sky130_fd_sc_hd__and4_1 _13464_ (.A(_01252_),
    .B(_05969_),
    .C(_02735_),
    .D(_02731_),
    .X(_05997_));
 sky130_fd_sc_hd__nor2_1 _13465_ (.A(_05996_),
    .B(_05997_),
    .Y(_05998_));
 sky130_fd_sc_hd__nand2_1 _13466_ (.A(_05985_),
    .B(_02722_),
    .Y(_06000_));
 sky130_fd_sc_hd__xnor2_1 _13467_ (.A(_05998_),
    .B(_06000_),
    .Y(_06001_));
 sky130_fd_sc_hd__nand2_1 _13468_ (.A(_05994_),
    .B(_06001_),
    .Y(_06002_));
 sky130_fd_sc_hd__or2_1 _13469_ (.A(_05994_),
    .B(_06001_),
    .X(_06003_));
 sky130_fd_sc_hd__nand2_1 _13470_ (.A(_06002_),
    .B(_06003_),
    .Y(_06004_));
 sky130_fd_sc_hd__a21oi_1 _13471_ (.A1(_05993_),
    .A2(_05989_),
    .B1(_06004_),
    .Y(_06005_));
 sky130_fd_sc_hd__and3_1 _13472_ (.A(_05993_),
    .B(_05989_),
    .C(_06004_),
    .X(_06006_));
 sky130_fd_sc_hd__nor2_1 _13473_ (.A(_06005_),
    .B(_06006_),
    .Y(_06007_));
 sky130_fd_sc_hd__xnor2_1 _13474_ (.A(_05992_),
    .B(_06007_),
    .Y(_06008_));
 sky130_fd_sc_hd__buf_2 _13475_ (.A(_02856_),
    .X(_06009_));
 sky130_fd_sc_hd__and4_1 _13476_ (.A(_01414_),
    .B(_06009_),
    .C(_01956_),
    .D(_03687_),
    .X(_06011_));
 sky130_fd_sc_hd__a22o_1 _13477_ (.A1(_06009_),
    .A2(_01956_),
    .B1(_03687_),
    .B2(_01414_),
    .X(_06012_));
 sky130_fd_sc_hd__and4b_1 _13478_ (.A_N(_06011_),
    .B(_06012_),
    .C(_01062_),
    .D(_03684_),
    .X(_06013_));
 sky130_fd_sc_hd__inv_2 _13479_ (.A(_06012_),
    .Y(_06014_));
 sky130_fd_sc_hd__o2bb2a_1 _13480_ (.A1_N(_01108_),
    .A2_N(_03697_),
    .B1(_06011_),
    .B2(_06014_),
    .X(_06015_));
 sky130_fd_sc_hd__and4_1 _13481_ (.A(_01062_),
    .B(_01415_),
    .C(_01958_),
    .D(_03690_),
    .X(_06016_));
 sky130_fd_sc_hd__or3b_1 _13482_ (.A(_06013_),
    .B(_06015_),
    .C_N(_06016_),
    .X(_06017_));
 sky130_fd_sc_hd__buf_2 _13483_ (.A(_02858_),
    .X(_06018_));
 sky130_fd_sc_hd__and4_1 _13484_ (.A(_06009_),
    .B(_06018_),
    .C(_01957_),
    .D(_03690_),
    .X(_06019_));
 sky130_fd_sc_hd__a22o_1 _13485_ (.A1(_06018_),
    .A2(_01957_),
    .B1(_03690_),
    .B2(_06009_),
    .X(_06020_));
 sky130_fd_sc_hd__and2b_1 _13486_ (.A_N(_06019_),
    .B(_06020_),
    .X(_06022_));
 sky130_fd_sc_hd__nand2_1 _13487_ (.A(_01415_),
    .B(_03697_),
    .Y(_06023_));
 sky130_fd_sc_hd__xnor2_1 _13488_ (.A(_06022_),
    .B(_06023_),
    .Y(_06024_));
 sky130_fd_sc_hd__o211ai_2 _13489_ (.A1(_06011_),
    .A2(_06013_),
    .B1(_01062_),
    .C1(_03699_),
    .Y(_06025_));
 sky130_fd_sc_hd__a211o_1 _13490_ (.A1(_01062_),
    .A2(_03699_),
    .B1(_06011_),
    .C1(_06013_),
    .X(_06026_));
 sky130_fd_sc_hd__and2_1 _13491_ (.A(_06025_),
    .B(_06026_),
    .X(_06027_));
 sky130_fd_sc_hd__nand2_1 _13492_ (.A(_06024_),
    .B(_06027_),
    .Y(_06028_));
 sky130_fd_sc_hd__or2_1 _13493_ (.A(_06024_),
    .B(_06027_),
    .X(_06029_));
 sky130_fd_sc_hd__nand2_1 _13494_ (.A(_06028_),
    .B(_06029_),
    .Y(_06030_));
 sky130_fd_sc_hd__nor2_1 _13495_ (.A(_06017_),
    .B(_06030_),
    .Y(_06031_));
 sky130_fd_sc_hd__a31o_1 _13496_ (.A1(_01415_),
    .A2(_03697_),
    .A3(_06020_),
    .B1(_06019_),
    .X(_06033_));
 sky130_fd_sc_hd__nand2_1 _13497_ (.A(_06009_),
    .B(_03684_),
    .Y(_06034_));
 sky130_fd_sc_hd__a21boi_1 _13498_ (.A1(_06018_),
    .A2(_03690_),
    .B1_N(_06034_),
    .Y(_06035_));
 sky130_fd_sc_hd__and4_1 _13499_ (.A(_06009_),
    .B(_06018_),
    .C(_03687_),
    .D(_03684_),
    .X(_06036_));
 sky130_fd_sc_hd__and4bb_1 _13500_ (.A_N(_06035_),
    .B_N(_06036_),
    .C(_01415_),
    .D(_03680_),
    .X(_06037_));
 sky130_fd_sc_hd__o2bb2a_1 _13501_ (.A1_N(_01415_),
    .A2_N(_03680_),
    .B1(_06035_),
    .B2(_06036_),
    .X(_06038_));
 sky130_fd_sc_hd__nor2_1 _13502_ (.A(_06037_),
    .B(_06038_),
    .Y(_06039_));
 sky130_fd_sc_hd__nand2_1 _13503_ (.A(_06033_),
    .B(_06039_),
    .Y(_06040_));
 sky130_fd_sc_hd__or2_1 _13504_ (.A(_06033_),
    .B(_06039_),
    .X(_06041_));
 sky130_fd_sc_hd__nand2_1 _13505_ (.A(_06040_),
    .B(_06041_),
    .Y(_06042_));
 sky130_fd_sc_hd__a21oi_1 _13506_ (.A1(_06025_),
    .A2(_06028_),
    .B1(_06042_),
    .Y(_06044_));
 sky130_fd_sc_hd__and3_1 _13507_ (.A(_06025_),
    .B(_06028_),
    .C(_06042_),
    .X(_06045_));
 sky130_fd_sc_hd__nor2_1 _13508_ (.A(_06044_),
    .B(_06045_),
    .Y(_06046_));
 sky130_fd_sc_hd__xnor2_1 _13509_ (.A(_06031_),
    .B(_06046_),
    .Y(_06047_));
 sky130_fd_sc_hd__nor2_2 _13510_ (.A(_06008_),
    .B(_06047_),
    .Y(_06048_));
 sky130_fd_sc_hd__a31o_1 _13511_ (.A1(_05985_),
    .A2(_02722_),
    .A3(_05998_),
    .B1(_05997_),
    .X(_06049_));
 sky130_fd_sc_hd__a22o_1 _13512_ (.A1(_05985_),
    .A2(_02736_),
    .B1(_02737_),
    .B2(_05969_),
    .X(_06050_));
 sky130_fd_sc_hd__nand4_1 _13513_ (.A(_05969_),
    .B(_05985_),
    .C(_02736_),
    .D(_02737_),
    .Y(_06051_));
 sky130_fd_sc_hd__nand2_1 _13514_ (.A(_06050_),
    .B(_06051_),
    .Y(_06052_));
 sky130_fd_sc_hd__xnor2_1 _13515_ (.A(_06049_),
    .B(_06052_),
    .Y(_06053_));
 sky130_fd_sc_hd__xor2_1 _13516_ (.A(_06002_),
    .B(_06053_),
    .X(_06055_));
 sky130_fd_sc_hd__a21oi_1 _13517_ (.A1(_05992_),
    .A2(_06007_),
    .B1(_06005_),
    .Y(_06056_));
 sky130_fd_sc_hd__nor2_1 _13518_ (.A(_06055_),
    .B(_06056_),
    .Y(_06057_));
 sky130_fd_sc_hd__and2_1 _13519_ (.A(_06055_),
    .B(_06056_),
    .X(_06058_));
 sky130_fd_sc_hd__nor2_1 _13520_ (.A(_06057_),
    .B(_06058_),
    .Y(_06059_));
 sky130_fd_sc_hd__a22o_1 _13521_ (.A1(_06018_),
    .A2(_03697_),
    .B1(_03699_),
    .B2(_06009_),
    .X(_06060_));
 sky130_fd_sc_hd__nand4_1 _13522_ (.A(_06009_),
    .B(_06018_),
    .C(_03697_),
    .D(_03699_),
    .Y(_06061_));
 sky130_fd_sc_hd__o211a_1 _13523_ (.A1(_06036_),
    .A2(_06037_),
    .B1(_06060_),
    .C1(_06061_),
    .X(_06062_));
 sky130_fd_sc_hd__a211oi_1 _13524_ (.A1(_06060_),
    .A2(_06061_),
    .B1(_06036_),
    .C1(_06037_),
    .Y(_06063_));
 sky130_fd_sc_hd__nor2_1 _13525_ (.A(_06062_),
    .B(_06063_),
    .Y(_06064_));
 sky130_fd_sc_hd__xor2_1 _13526_ (.A(_06040_),
    .B(_06064_),
    .X(_06066_));
 sky130_fd_sc_hd__a21oi_1 _13527_ (.A1(_06031_),
    .A2(_06046_),
    .B1(_06044_),
    .Y(_06067_));
 sky130_fd_sc_hd__nor2_1 _13528_ (.A(_06066_),
    .B(_06067_),
    .Y(_06068_));
 sky130_fd_sc_hd__and2_1 _13529_ (.A(_06066_),
    .B(_06067_),
    .X(_06069_));
 sky130_fd_sc_hd__nor2_1 _13530_ (.A(_06068_),
    .B(_06069_),
    .Y(_06070_));
 sky130_fd_sc_hd__nand2_1 _13531_ (.A(_06059_),
    .B(_06070_),
    .Y(_06071_));
 sky130_fd_sc_hd__or2_1 _13532_ (.A(_06059_),
    .B(_06070_),
    .X(_06072_));
 sky130_fd_sc_hd__and2_1 _13533_ (.A(_06071_),
    .B(_06072_),
    .X(_06073_));
 sky130_fd_sc_hd__buf_2 _13534_ (.A(_02766_),
    .X(_06074_));
 sky130_fd_sc_hd__buf_2 _13535_ (.A(_01958_),
    .X(_06075_));
 sky130_fd_sc_hd__buf_2 _13536_ (.A(_02722_),
    .X(_06077_));
 sky130_fd_sc_hd__buf_2 _13537_ (.A(_03690_),
    .X(_06078_));
 sky130_fd_sc_hd__and4_1 _13538_ (.A(_06074_),
    .B(_06075_),
    .C(_06077_),
    .D(_06078_),
    .X(_06079_));
 sky130_fd_sc_hd__a22oi_1 _13539_ (.A1(_06075_),
    .A2(_06077_),
    .B1(_06078_),
    .B2(_06074_),
    .Y(_06080_));
 sky130_fd_sc_hd__nor2_1 _13540_ (.A(_06079_),
    .B(_06080_),
    .Y(_06081_));
 sky130_fd_sc_hd__a21oi_1 _13541_ (.A1(_06048_),
    .A2(_06073_),
    .B1(_06081_),
    .Y(_06082_));
 sky130_fd_sc_hd__o21ba_1 _13542_ (.A1(_06048_),
    .A2(_06073_),
    .B1_N(_06082_),
    .X(_06083_));
 sky130_fd_sc_hd__and3_1 _13543_ (.A(_05994_),
    .B(_06001_),
    .C(_06053_),
    .X(_06084_));
 sky130_fd_sc_hd__and3_1 _13544_ (.A(_06049_),
    .B(_06050_),
    .C(_06051_),
    .X(_06085_));
 sky130_fd_sc_hd__and3_1 _13545_ (.A(_05985_),
    .B(_02737_),
    .C(_05995_),
    .X(_06086_));
 sky130_fd_sc_hd__xor2_1 _13546_ (.A(_06085_),
    .B(_06086_),
    .X(_06088_));
 sky130_fd_sc_hd__nor3_1 _13547_ (.A(_06084_),
    .B(_06057_),
    .C(_06088_),
    .Y(_06089_));
 sky130_fd_sc_hd__o21a_1 _13548_ (.A1(_06084_),
    .A2(_06057_),
    .B1(_06088_),
    .X(_06090_));
 sky130_fd_sc_hd__nor2_1 _13549_ (.A(_06089_),
    .B(_06090_),
    .Y(_06091_));
 sky130_fd_sc_hd__and3_1 _13550_ (.A(_06033_),
    .B(_06039_),
    .C(_06064_),
    .X(_06092_));
 sky130_fd_sc_hd__and3_1 _13551_ (.A(_06018_),
    .B(_04013_),
    .C(_06034_),
    .X(_06093_));
 sky130_fd_sc_hd__xor2_1 _13552_ (.A(_06062_),
    .B(_06093_),
    .X(_06094_));
 sky130_fd_sc_hd__nor3_1 _13553_ (.A(_06092_),
    .B(_06068_),
    .C(_06094_),
    .Y(_06095_));
 sky130_fd_sc_hd__o21a_1 _13554_ (.A1(_06092_),
    .A2(_06068_),
    .B1(_06094_),
    .X(_06096_));
 sky130_fd_sc_hd__nor2_1 _13555_ (.A(_06095_),
    .B(_06096_),
    .Y(_06097_));
 sky130_fd_sc_hd__nand2_1 _13556_ (.A(_06091_),
    .B(_06097_),
    .Y(_06099_));
 sky130_fd_sc_hd__or2_1 _13557_ (.A(_06091_),
    .B(_06097_),
    .X(_06100_));
 sky130_fd_sc_hd__nand2_1 _13558_ (.A(_06099_),
    .B(_06100_),
    .Y(_06101_));
 sky130_fd_sc_hd__and2_1 _13559_ (.A(_06071_),
    .B(_06101_),
    .X(_06102_));
 sky130_fd_sc_hd__nor2_1 _13560_ (.A(_06071_),
    .B(_06101_),
    .Y(_06103_));
 sky130_fd_sc_hd__a22o_1 _13561_ (.A1(_06077_),
    .A2(_06078_),
    .B1(_02736_),
    .B2(_01958_),
    .X(_06104_));
 sky130_fd_sc_hd__nand4_1 _13562_ (.A(_06075_),
    .B(_06077_),
    .C(_06078_),
    .D(_02736_),
    .Y(_06105_));
 sky130_fd_sc_hd__a22oi_1 _13563_ (.A1(_06074_),
    .A2(_04014_),
    .B1(_06104_),
    .B2(_06105_),
    .Y(_06106_));
 sky130_fd_sc_hd__and4_1 _13564_ (.A(_06074_),
    .B(_04014_),
    .C(_06104_),
    .D(_06105_),
    .X(_06107_));
 sky130_fd_sc_hd__or2_1 _13565_ (.A(_06106_),
    .B(_06107_),
    .X(_06108_));
 sky130_fd_sc_hd__xnor2_1 _13566_ (.A(_06108_),
    .B(_06079_),
    .Y(_06110_));
 sky130_fd_sc_hd__or2_1 _13567_ (.A(_06103_),
    .B(_06110_),
    .X(_06111_));
 sky130_fd_sc_hd__o21ai_1 _13568_ (.A1(_06102_),
    .A2(_06103_),
    .B1(_06110_),
    .Y(_06112_));
 sky130_fd_sc_hd__o21a_1 _13569_ (.A1(_06102_),
    .A2(_06111_),
    .B1(_06112_),
    .X(_06113_));
 sky130_fd_sc_hd__and2b_1 _13570_ (.A_N(_06083_),
    .B(_06113_),
    .X(_06114_));
 sky130_fd_sc_hd__and2b_1 _13571_ (.A_N(_06113_),
    .B(_06083_),
    .X(_06115_));
 sky130_fd_sc_hd__nor2_2 _13572_ (.A(_06114_),
    .B(_06115_),
    .Y(_06116_));
 sky130_fd_sc_hd__and2_1 _13573_ (.A(_05978_),
    .B(_05991_),
    .X(_06117_));
 sky130_fd_sc_hd__nor2_1 _13574_ (.A(_05992_),
    .B(_06117_),
    .Y(_06118_));
 sky130_fd_sc_hd__and4_1 _13575_ (.A(_06009_),
    .B(_05969_),
    .C(_06018_),
    .D(_05985_),
    .X(_06119_));
 sky130_fd_sc_hd__nand2_1 _13576_ (.A(_02855_),
    .B(_03785_),
    .Y(_06121_));
 sky130_fd_sc_hd__and4_1 _13577_ (.A(_01249_),
    .B(_02855_),
    .C(_03785_),
    .D(_02857_),
    .X(_06122_));
 sky130_fd_sc_hd__a21boi_1 _13578_ (.A1(_01250_),
    .A2(_02858_),
    .B1_N(_06121_),
    .Y(_06123_));
 sky130_fd_sc_hd__nor2_1 _13579_ (.A(_06122_),
    .B(_06123_),
    .Y(_06124_));
 sky130_fd_sc_hd__and3_1 _13580_ (.A(_01414_),
    .B(_03783_),
    .C(_06124_),
    .X(_06125_));
 sky130_fd_sc_hd__or2_1 _13581_ (.A(_06122_),
    .B(_06125_),
    .X(_06126_));
 sky130_fd_sc_hd__nand4_1 _13582_ (.A(_06009_),
    .B(_03785_),
    .C(_02858_),
    .D(_03783_),
    .Y(_06127_));
 sky130_fd_sc_hd__a22o_1 _13583_ (.A1(_03785_),
    .A2(_02858_),
    .B1(_03783_),
    .B2(_02856_),
    .X(_06128_));
 sky130_fd_sc_hd__and3_1 _13584_ (.A(_06126_),
    .B(_06127_),
    .C(_06128_),
    .X(_06129_));
 sky130_fd_sc_hd__and4_1 _13585_ (.A(_06018_),
    .B(_05985_),
    .C(_06121_),
    .D(_06129_),
    .X(_06130_));
 sky130_fd_sc_hd__a31o_1 _13586_ (.A1(_06018_),
    .A2(_05985_),
    .A3(_06121_),
    .B1(_06129_),
    .X(_06132_));
 sky130_fd_sc_hd__and2b_1 _13587_ (.A_N(_06130_),
    .B(_06132_),
    .X(_06133_));
 sky130_fd_sc_hd__a21oi_1 _13588_ (.A1(_01414_),
    .A2(_03783_),
    .B1(_06124_),
    .Y(_06134_));
 sky130_fd_sc_hd__or2_1 _13589_ (.A(_06125_),
    .B(_06134_),
    .X(_06135_));
 sky130_fd_sc_hd__and4_1 _13590_ (.A(_01181_),
    .B(_01250_),
    .C(_02856_),
    .D(_02858_),
    .X(_06136_));
 sky130_fd_sc_hd__a22oi_1 _13591_ (.A1(_01250_),
    .A2(_02856_),
    .B1(_02858_),
    .B2(_01181_),
    .Y(_06137_));
 sky130_fd_sc_hd__and4bb_1 _13592_ (.A_N(_06136_),
    .B_N(_06137_),
    .C(_01414_),
    .D(_03785_),
    .X(_06138_));
 sky130_fd_sc_hd__or2_1 _13593_ (.A(_06136_),
    .B(_06138_),
    .X(_06139_));
 sky130_fd_sc_hd__and2b_1 _13594_ (.A_N(_06135_),
    .B(_06139_),
    .X(_06140_));
 sky130_fd_sc_hd__a21oi_1 _13595_ (.A1(_06127_),
    .A2(_06128_),
    .B1(_06126_),
    .Y(_06141_));
 sky130_fd_sc_hd__nor2_1 _13596_ (.A(_06129_),
    .B(_06141_),
    .Y(_06143_));
 sky130_fd_sc_hd__a22o_1 _13597_ (.A1(_01413_),
    .A2(_01249_),
    .B1(_02856_),
    .B2(_01180_),
    .X(_06144_));
 sky130_fd_sc_hd__and3_1 _13598_ (.A(_01181_),
    .B(_01413_),
    .C(_01250_),
    .X(_06145_));
 sky130_fd_sc_hd__a32o_1 _13599_ (.A1(_01061_),
    .A2(_03785_),
    .A3(_06144_),
    .B1(_06145_),
    .B2(_02856_),
    .X(_06146_));
 sky130_fd_sc_hd__and3_1 _13600_ (.A(_01061_),
    .B(_03783_),
    .C(_06146_),
    .X(_06147_));
 sky130_fd_sc_hd__o2bb2a_1 _13601_ (.A1_N(_01414_),
    .A2_N(_03785_),
    .B1(_06136_),
    .B2(_06137_),
    .X(_06148_));
 sky130_fd_sc_hd__a21oi_1 _13602_ (.A1(_01061_),
    .A2(_03783_),
    .B1(_06146_),
    .Y(_06149_));
 sky130_fd_sc_hd__nor4_1 _13603_ (.A(_06138_),
    .B(_06147_),
    .C(_06148_),
    .D(_06149_),
    .Y(_06150_));
 sky130_fd_sc_hd__xnor2_1 _13604_ (.A(_06139_),
    .B(_06135_),
    .Y(_06151_));
 sky130_fd_sc_hd__o21a_1 _13605_ (.A1(_06147_),
    .A2(net141),
    .B1(_06151_),
    .X(_06152_));
 sky130_fd_sc_hd__a21bo_1 _13606_ (.A1(_02856_),
    .A2(_06145_),
    .B1_N(_06144_),
    .X(_06154_));
 sky130_fd_sc_hd__nand2_1 _13607_ (.A(_01061_),
    .B(_03785_),
    .Y(_06155_));
 sky130_fd_sc_hd__xnor2_1 _13608_ (.A(_06154_),
    .B(_06155_),
    .Y(_06156_));
 sky130_fd_sc_hd__nor2_1 _13609_ (.A(_05951_),
    .B(_06156_),
    .Y(_06157_));
 sky130_fd_sc_hd__o22a_1 _13610_ (.A1(_06138_),
    .A2(_06148_),
    .B1(_06149_),
    .B2(_06147_),
    .X(_06158_));
 sky130_fd_sc_hd__nor2_1 _13611_ (.A(_06150_),
    .B(_06158_),
    .Y(_06159_));
 sky130_fd_sc_hd__nand2_1 _13612_ (.A(_06157_),
    .B(_06159_),
    .Y(_06160_));
 sky130_fd_sc_hd__nor3_1 _13613_ (.A(_06147_),
    .B(net141),
    .C(_06151_),
    .Y(_06161_));
 sky130_fd_sc_hd__or3_1 _13614_ (.A(_06152_),
    .B(_06160_),
    .C(_06161_),
    .X(_06162_));
 sky130_fd_sc_hd__and2b_1 _13615_ (.A_N(_06152_),
    .B(_06162_),
    .X(_06163_));
 sky130_fd_sc_hd__xor2_1 _13616_ (.A(_06140_),
    .B(_06143_),
    .X(_06165_));
 sky130_fd_sc_hd__and2b_1 _13617_ (.A_N(_06163_),
    .B(_06165_),
    .X(_06166_));
 sky130_fd_sc_hd__a21o_1 _13618_ (.A1(_06140_),
    .A2(_06143_),
    .B1(_06166_),
    .X(_06167_));
 sky130_fd_sc_hd__and2_1 _13619_ (.A(_06133_),
    .B(_06167_),
    .X(_06168_));
 sky130_fd_sc_hd__or4_1 _13620_ (.A(_06118_),
    .B(_06119_),
    .C(_06130_),
    .D(_06168_),
    .X(_06169_));
 sky130_fd_sc_hd__o31ai_1 _13621_ (.A1(_06119_),
    .A2(_06130_),
    .A3(_06168_),
    .B1(_06118_),
    .Y(_06170_));
 sky130_fd_sc_hd__and2_1 _13622_ (.A(_06017_),
    .B(_06030_),
    .X(_06171_));
 sky130_fd_sc_hd__or2_1 _13623_ (.A(_06031_),
    .B(_06171_),
    .X(_06172_));
 sky130_fd_sc_hd__nand2_1 _13624_ (.A(_06170_),
    .B(_06172_),
    .Y(_06173_));
 sky130_fd_sc_hd__and2_1 _13625_ (.A(_06008_),
    .B(_06047_),
    .X(_06174_));
 sky130_fd_sc_hd__nor2_1 _13626_ (.A(_06048_),
    .B(_06174_),
    .Y(_06176_));
 sky130_fd_sc_hd__a21oi_1 _13627_ (.A1(_06169_),
    .A2(_06173_),
    .B1(_06176_),
    .Y(_06177_));
 sky130_fd_sc_hd__and3_1 _13628_ (.A(_06176_),
    .B(_06169_),
    .C(_06173_),
    .X(_06178_));
 sky130_fd_sc_hd__a21oi_1 _13629_ (.A1(_06074_),
    .A2(_06075_),
    .B1(_06178_),
    .Y(_06179_));
 sky130_fd_sc_hd__or2_1 _13630_ (.A(_06177_),
    .B(_06179_),
    .X(_06180_));
 sky130_fd_sc_hd__or2_1 _13631_ (.A(_06048_),
    .B(_06073_),
    .X(_06181_));
 sky130_fd_sc_hd__nand2_1 _13632_ (.A(_06048_),
    .B(_06073_),
    .Y(_06182_));
 sky130_fd_sc_hd__nand2_1 _13633_ (.A(_06181_),
    .B(_06182_),
    .Y(_06183_));
 sky130_fd_sc_hd__a22o_1 _13634_ (.A1(_06181_),
    .A2(_06082_),
    .B1(_06183_),
    .B2(_06081_),
    .X(_06184_));
 sky130_fd_sc_hd__and2b_1 _13635_ (.A_N(_06180_),
    .B(_06184_),
    .X(_06185_));
 sky130_fd_sc_hd__and2b_1 _13636_ (.A_N(_06184_),
    .B(_06180_),
    .X(_06187_));
 sky130_fd_sc_hd__nor2_1 _13637_ (.A(_06185_),
    .B(_06187_),
    .Y(_06188_));
 sky130_fd_sc_hd__inv_2 _13638_ (.A(_06188_),
    .Y(_06189_));
 sky130_fd_sc_hd__nand2_1 _13639_ (.A(_06169_),
    .B(_06170_),
    .Y(_06190_));
 sky130_fd_sc_hd__xor2_1 _13640_ (.A(_06172_),
    .B(_06190_),
    .X(_06191_));
 sky130_fd_sc_hd__or2_1 _13641_ (.A(_05975_),
    .B(_05976_),
    .X(_06192_));
 sky130_fd_sc_hd__nand2_1 _13642_ (.A(_05978_),
    .B(_06192_),
    .Y(_06193_));
 sky130_fd_sc_hd__xnor2_1 _13643_ (.A(_06133_),
    .B(_06167_),
    .Y(_06194_));
 sky130_fd_sc_hd__nand2_1 _13644_ (.A(_06193_),
    .B(_06194_),
    .Y(_06195_));
 sky130_fd_sc_hd__nor2_1 _13645_ (.A(_06193_),
    .B(_06194_),
    .Y(_06196_));
 sky130_fd_sc_hd__or2_1 _13646_ (.A(_06013_),
    .B(_06015_),
    .X(_06198_));
 sky130_fd_sc_hd__xnor2_1 _13647_ (.A(_06198_),
    .B(_06016_),
    .Y(_06199_));
 sky130_fd_sc_hd__or2_1 _13648_ (.A(_06196_),
    .B(_06199_),
    .X(_06200_));
 sky130_fd_sc_hd__and3_1 _13649_ (.A(_06191_),
    .B(_06195_),
    .C(_06200_),
    .X(_06201_));
 sky130_fd_sc_hd__a21oi_1 _13650_ (.A1(_06195_),
    .A2(_06200_),
    .B1(_06191_),
    .Y(_06202_));
 sky130_fd_sc_hd__or2_1 _13651_ (.A(_06201_),
    .B(_06202_),
    .X(_06203_));
 sky130_fd_sc_hd__inv_2 _13652_ (.A(_06195_),
    .Y(_06204_));
 sky130_fd_sc_hd__nor2_1 _13653_ (.A(_06204_),
    .B(_06196_),
    .Y(_06205_));
 sky130_fd_sc_hd__xnor2_1 _13654_ (.A(_06199_),
    .B(_06205_),
    .Y(_06206_));
 sky130_fd_sc_hd__inv_2 _13655_ (.A(_05976_),
    .Y(_06207_));
 sky130_fd_sc_hd__a22o_1 _13656_ (.A1(_01252_),
    .A2(_02766_),
    .B1(_06077_),
    .B2(_01183_),
    .X(_06209_));
 sky130_fd_sc_hd__and2b_1 _13657_ (.A_N(_06165_),
    .B(_06163_),
    .X(_06210_));
 sky130_fd_sc_hd__nor2_1 _13658_ (.A(_06166_),
    .B(_06210_),
    .Y(_06211_));
 sky130_fd_sc_hd__a21o_1 _13659_ (.A1(_06207_),
    .A2(_06209_),
    .B1(_06211_),
    .X(_06212_));
 sky130_fd_sc_hd__a22oi_1 _13660_ (.A1(_01415_),
    .A2(_01958_),
    .B1(_06078_),
    .B2(_01108_),
    .Y(_06213_));
 sky130_fd_sc_hd__nor2_1 _13661_ (.A(_06016_),
    .B(_06213_),
    .Y(_06214_));
 sky130_fd_sc_hd__nand3_1 _13662_ (.A(_06207_),
    .B(_06209_),
    .C(_06211_),
    .Y(_06215_));
 sky130_fd_sc_hd__a21bo_1 _13663_ (.A1(_06212_),
    .A2(_06214_),
    .B1_N(_06215_),
    .X(_06216_));
 sky130_fd_sc_hd__or2b_1 _13664_ (.A(_06206_),
    .B_N(_06216_),
    .X(_06217_));
 sky130_fd_sc_hd__or2b_1 _13665_ (.A(_06216_),
    .B_N(_06206_),
    .X(_06218_));
 sky130_fd_sc_hd__nand2_2 _13666_ (.A(_06217_),
    .B(_06218_),
    .Y(_06220_));
 sky130_fd_sc_hd__nand2_1 _13667_ (.A(_01108_),
    .B(_06075_),
    .Y(_06221_));
 sky130_fd_sc_hd__o21ai_1 _13668_ (.A1(_06152_),
    .A2(_06161_),
    .B1(_06160_),
    .Y(_06222_));
 sky130_fd_sc_hd__and2_1 _13669_ (.A(_06162_),
    .B(_06222_),
    .X(_06223_));
 sky130_fd_sc_hd__nand3_1 _13670_ (.A(_01183_),
    .B(_06074_),
    .C(_06223_),
    .Y(_06224_));
 sky130_fd_sc_hd__a21oi_1 _13671_ (.A1(_01183_),
    .A2(_02766_),
    .B1(_06223_),
    .Y(_06225_));
 sky130_fd_sc_hd__a21o_1 _13672_ (.A1(_06221_),
    .A2(_06224_),
    .B1(_06225_),
    .X(_06226_));
 sky130_fd_sc_hd__nand2_1 _13673_ (.A(_06215_),
    .B(_06212_),
    .Y(_06227_));
 sky130_fd_sc_hd__xor2_2 _13674_ (.A(_06214_),
    .B(_06227_),
    .X(_06228_));
 sky130_fd_sc_hd__o31a_1 _13675_ (.A1(_06220_),
    .A2(_06226_),
    .A3(_06228_),
    .B1(_06217_),
    .X(_06229_));
 sky130_fd_sc_hd__nor2_1 _13676_ (.A(_06203_),
    .B(_06229_),
    .Y(_06231_));
 sky130_fd_sc_hd__o211ai_1 _13677_ (.A1(_06177_),
    .A2(_06178_),
    .B1(_06074_),
    .C1(_06075_),
    .Y(_06232_));
 sky130_fd_sc_hd__a211o_1 _13678_ (.A1(_06074_),
    .A2(_06075_),
    .B1(_06177_),
    .C1(_06178_),
    .X(_06233_));
 sky130_fd_sc_hd__nand2_1 _13679_ (.A(_06232_),
    .B(_06233_),
    .Y(_06234_));
 sky130_fd_sc_hd__o21ai_1 _13680_ (.A1(_06201_),
    .A2(_06231_),
    .B1(_06234_),
    .Y(_06235_));
 sky130_fd_sc_hd__nor2_1 _13681_ (.A(_06189_),
    .B(_06235_),
    .Y(_06236_));
 sky130_fd_sc_hd__or2_2 _13682_ (.A(_06185_),
    .B(_06236_),
    .X(_06237_));
 sky130_fd_sc_hd__xnor2_4 _13683_ (.A(_06116_),
    .B(_06237_),
    .Y(_06238_));
 sky130_fd_sc_hd__and2_1 _13684_ (.A(_06189_),
    .B(_06235_),
    .X(_06239_));
 sky130_fd_sc_hd__or2_1 _13685_ (.A(_06236_),
    .B(_06239_),
    .X(_06240_));
 sky130_fd_sc_hd__and4_1 _13686_ (.A(_02427_),
    .B(_02426_),
    .C(_02735_),
    .D(_02731_),
    .X(_06242_));
 sky130_fd_sc_hd__and4_1 _13687_ (.A(_01288_),
    .B(_02090_),
    .C(_02725_),
    .D(_02728_),
    .X(_06243_));
 sky130_fd_sc_hd__nand2_1 _13688_ (.A(_02090_),
    .B(_02725_),
    .Y(_06244_));
 sky130_fd_sc_hd__a21boi_1 _13689_ (.A1(_01289_),
    .A2(_02730_),
    .B1_N(_06244_),
    .Y(_06245_));
 sky130_fd_sc_hd__nor2_1 _13690_ (.A(_06243_),
    .B(_06245_),
    .Y(_06246_));
 sky130_fd_sc_hd__and3_1 _13691_ (.A(_02088_),
    .B(_02720_),
    .C(_06246_),
    .X(_06247_));
 sky130_fd_sc_hd__a22oi_1 _13692_ (.A1(_02426_),
    .A2(_02736_),
    .B1(_02737_),
    .B2(_02427_),
    .Y(_06248_));
 sky130_fd_sc_hd__nor2_1 _13693_ (.A(_06242_),
    .B(_06248_),
    .Y(_06249_));
 sky130_fd_sc_hd__o21a_1 _13694_ (.A1(_06243_),
    .A2(_06247_),
    .B1(_06249_),
    .X(_06250_));
 sky130_fd_sc_hd__and3_1 _13695_ (.A(_02426_),
    .B(_02737_),
    .C(_06244_),
    .X(_06251_));
 sky130_fd_sc_hd__and2_1 _13696_ (.A(_06250_),
    .B(_06251_),
    .X(_06253_));
 sky130_fd_sc_hd__and4_1 _13697_ (.A(_00416_),
    .B(_01288_),
    .C(_02725_),
    .D(_02730_),
    .X(_06254_));
 sky130_fd_sc_hd__a22oi_1 _13698_ (.A1(_01289_),
    .A2(_02726_),
    .B1(_02730_),
    .B2(_01188_),
    .Y(_06255_));
 sky130_fd_sc_hd__and4bb_1 _13699_ (.A_N(_06254_),
    .B_N(_06255_),
    .C(_02427_),
    .D(_02720_),
    .X(_06256_));
 sky130_fd_sc_hd__nor2_1 _13700_ (.A(_06254_),
    .B(_06256_),
    .Y(_06257_));
 sky130_fd_sc_hd__a21oi_1 _13701_ (.A1(_02426_),
    .A2(_02721_),
    .B1(_06246_),
    .Y(_06258_));
 sky130_fd_sc_hd__or3_1 _13702_ (.A(_06247_),
    .B(_06257_),
    .C(_06258_),
    .X(_06259_));
 sky130_fd_sc_hd__nor3_1 _13703_ (.A(_06243_),
    .B(_06247_),
    .C(_06249_),
    .Y(_06260_));
 sky130_fd_sc_hd__nor2_1 _13704_ (.A(_06250_),
    .B(_06260_),
    .Y(_06261_));
 sky130_fd_sc_hd__and2b_1 _13705_ (.A_N(_06259_),
    .B(_06261_),
    .X(_06262_));
 sky130_fd_sc_hd__a22o_1 _13706_ (.A1(_01288_),
    .A2(_02720_),
    .B1(_02725_),
    .B2(_00416_),
    .X(_06264_));
 sky130_fd_sc_hd__a21bo_1 _13707_ (.A1(_02726_),
    .A2(_05887_),
    .B1_N(_06264_),
    .X(_06265_));
 sky130_fd_sc_hd__nand2_1 _13708_ (.A(_02427_),
    .B(_02759_),
    .Y(_06266_));
 sky130_fd_sc_hd__xor2_1 _13709_ (.A(_06265_),
    .B(_06266_),
    .X(_06267_));
 sky130_fd_sc_hd__and3_1 _13710_ (.A(_02759_),
    .B(_05887_),
    .C(_06267_),
    .X(_06268_));
 sky130_fd_sc_hd__o2bb2a_1 _13711_ (.A1_N(_02427_),
    .A2_N(_02721_),
    .B1(_06254_),
    .B2(_06255_),
    .X(_06269_));
 sky130_fd_sc_hd__or2_1 _13712_ (.A(_06256_),
    .B(_06269_),
    .X(_06270_));
 sky130_fd_sc_hd__a32o_1 _13713_ (.A1(_02427_),
    .A2(_02758_),
    .A3(_06264_),
    .B1(_05887_),
    .B2(_02726_),
    .X(_06271_));
 sky130_fd_sc_hd__and3_1 _13714_ (.A(_02426_),
    .B(_02759_),
    .C(_06271_),
    .X(_06272_));
 sky130_fd_sc_hd__a21oi_1 _13715_ (.A1(_02426_),
    .A2(_02759_),
    .B1(_06271_),
    .Y(_06273_));
 sky130_fd_sc_hd__nor2_1 _13716_ (.A(_06272_),
    .B(_06273_),
    .Y(_06275_));
 sky130_fd_sc_hd__xnor2_1 _13717_ (.A(_06270_),
    .B(_06275_),
    .Y(_06276_));
 sky130_fd_sc_hd__nand2_1 _13718_ (.A(_06268_),
    .B(_06276_),
    .Y(_06277_));
 sky130_fd_sc_hd__and2b_1 _13719_ (.A_N(_06270_),
    .B(_06275_),
    .X(_06278_));
 sky130_fd_sc_hd__o21ai_1 _13720_ (.A1(_06247_),
    .A2(_06258_),
    .B1(_06257_),
    .Y(_06279_));
 sky130_fd_sc_hd__and2_1 _13721_ (.A(_06259_),
    .B(_06279_),
    .X(_06280_));
 sky130_fd_sc_hd__o21ai_1 _13722_ (.A1(_06272_),
    .A2(_06278_),
    .B1(_06280_),
    .Y(_06281_));
 sky130_fd_sc_hd__or3_1 _13723_ (.A(_06272_),
    .B(_06278_),
    .C(_06280_),
    .X(_06282_));
 sky130_fd_sc_hd__nand2_1 _13724_ (.A(_06281_),
    .B(_06282_),
    .Y(_06283_));
 sky130_fd_sc_hd__o21a_1 _13725_ (.A1(_06277_),
    .A2(_06283_),
    .B1(_06281_),
    .X(_06284_));
 sky130_fd_sc_hd__xnor2_1 _13726_ (.A(_06259_),
    .B(_06261_),
    .Y(_06286_));
 sky130_fd_sc_hd__and2b_1 _13727_ (.A_N(_06284_),
    .B(_06286_),
    .X(_06287_));
 sky130_fd_sc_hd__nor2_1 _13728_ (.A(_06250_),
    .B(_06251_),
    .Y(_06288_));
 sky130_fd_sc_hd__nor2_1 _13729_ (.A(_06253_),
    .B(_06288_),
    .Y(_06289_));
 sky130_fd_sc_hd__o21a_1 _13730_ (.A1(_06262_),
    .A2(_06287_),
    .B1(_06289_),
    .X(_06290_));
 sky130_fd_sc_hd__and2b_1 _13731_ (.A_N(_06286_),
    .B(_06284_),
    .X(_06291_));
 sky130_fd_sc_hd__nor2_1 _13732_ (.A(_06287_),
    .B(_06291_),
    .Y(_06292_));
 sky130_fd_sc_hd__nor2_1 _13733_ (.A(_05855_),
    .B(_05859_),
    .Y(_06293_));
 sky130_fd_sc_hd__nand2_1 _13734_ (.A(_00915_),
    .B(_02725_),
    .Y(_06294_));
 sky130_fd_sc_hd__and3_1 _13735_ (.A(_00916_),
    .B(_02730_),
    .C(_06294_),
    .X(_06295_));
 sky130_fd_sc_hd__nand2_1 _13736_ (.A(_06293_),
    .B(_06295_),
    .Y(_06297_));
 sky130_fd_sc_hd__xor2_1 _13737_ (.A(_06293_),
    .B(_06295_),
    .X(_06298_));
 sky130_fd_sc_hd__o21ai_1 _13738_ (.A1(_05861_),
    .A2(_05866_),
    .B1(_06298_),
    .Y(_06299_));
 sky130_fd_sc_hd__and3_1 _13739_ (.A(_05858_),
    .B(_06297_),
    .C(_06299_),
    .X(_06300_));
 sky130_fd_sc_hd__nor2_1 _13740_ (.A(_05870_),
    .B(_05873_),
    .Y(_06301_));
 sky130_fd_sc_hd__nand2_1 _13741_ (.A(_02090_),
    .B(_02855_),
    .Y(_06302_));
 sky130_fd_sc_hd__and3_1 _13742_ (.A(_02088_),
    .B(_02858_),
    .C(_06302_),
    .X(_06303_));
 sky130_fd_sc_hd__xor2_1 _13743_ (.A(_06301_),
    .B(_06303_),
    .X(_06304_));
 sky130_fd_sc_hd__o21a_1 _13744_ (.A1(_05875_),
    .A2(_05881_),
    .B1(_06304_),
    .X(_06305_));
 sky130_fd_sc_hd__a21o_1 _13745_ (.A1(_06301_),
    .A2(_06303_),
    .B1(_06305_),
    .X(_06306_));
 sky130_fd_sc_hd__and2b_1 _13746_ (.A_N(_06306_),
    .B(_05872_),
    .X(_06308_));
 sky130_fd_sc_hd__nor2_1 _13747_ (.A(_06300_),
    .B(_06308_),
    .Y(_06309_));
 sky130_fd_sc_hd__xor2_1 _13748_ (.A(_06277_),
    .B(_06283_),
    .X(_06310_));
 sky130_fd_sc_hd__and3_1 _13749_ (.A(_06292_),
    .B(_06309_),
    .C(_06310_),
    .X(_06311_));
 sky130_fd_sc_hd__and2_1 _13750_ (.A(_06309_),
    .B(_06310_),
    .X(_06312_));
 sky130_fd_sc_hd__nor2_1 _13751_ (.A(_06309_),
    .B(_06310_),
    .Y(_06313_));
 sky130_fd_sc_hd__nor2_1 _13752_ (.A(_06312_),
    .B(_06313_),
    .Y(_06314_));
 sky130_fd_sc_hd__or3_1 _13753_ (.A(_05861_),
    .B(_05866_),
    .C(_06298_),
    .X(_06315_));
 sky130_fd_sc_hd__and2_1 _13754_ (.A(_06299_),
    .B(_06315_),
    .X(_06316_));
 sky130_fd_sc_hd__nor3_1 _13755_ (.A(_05875_),
    .B(_05881_),
    .C(_06304_),
    .Y(_06317_));
 sky130_fd_sc_hd__nor2_1 _13756_ (.A(_06305_),
    .B(_06317_),
    .Y(_06319_));
 sky130_fd_sc_hd__nand2_1 _13757_ (.A(_06316_),
    .B(_06319_),
    .Y(_06320_));
 sky130_fd_sc_hd__and2_1 _13758_ (.A(_06300_),
    .B(_06308_),
    .X(_06321_));
 sky130_fd_sc_hd__or2_1 _13759_ (.A(_06309_),
    .B(_06321_),
    .X(_06322_));
 sky130_fd_sc_hd__nand2_1 _13760_ (.A(_06320_),
    .B(_06322_),
    .Y(_06323_));
 sky130_fd_sc_hd__or2_1 _13761_ (.A(_06268_),
    .B(_06276_),
    .X(_06324_));
 sky130_fd_sc_hd__and2_1 _13762_ (.A(_06277_),
    .B(_06324_),
    .X(_06325_));
 sky130_fd_sc_hd__nor2_1 _13763_ (.A(_06320_),
    .B(_06322_),
    .Y(_06326_));
 sky130_fd_sc_hd__or2_1 _13764_ (.A(_06325_),
    .B(_06326_),
    .X(_06327_));
 sky130_fd_sc_hd__and3_1 _13765_ (.A(_06314_),
    .B(_06323_),
    .C(_06327_),
    .X(_06328_));
 sky130_fd_sc_hd__a21oi_1 _13766_ (.A1(_06323_),
    .A2(_06327_),
    .B1(_06314_),
    .Y(_06330_));
 sky130_fd_sc_hd__nor2_1 _13767_ (.A(_06328_),
    .B(_06330_),
    .Y(_06331_));
 sky130_fd_sc_hd__nand2_1 _13768_ (.A(_05867_),
    .B(_05882_),
    .Y(_06332_));
 sky130_fd_sc_hd__xnor2_1 _13769_ (.A(_06316_),
    .B(_06319_),
    .Y(_06333_));
 sky130_fd_sc_hd__and2_1 _13770_ (.A(_06332_),
    .B(_06333_),
    .X(_06334_));
 sky130_fd_sc_hd__inv_2 _13771_ (.A(_06334_),
    .Y(_06335_));
 sky130_fd_sc_hd__a21oi_1 _13772_ (.A1(_02765_),
    .A2(_05887_),
    .B1(_06267_),
    .Y(_06336_));
 sky130_fd_sc_hd__or2_1 _13773_ (.A(_06268_),
    .B(_06336_),
    .X(_06337_));
 sky130_fd_sc_hd__o21ai_1 _13774_ (.A1(_06332_),
    .A2(_06333_),
    .B1(_06337_),
    .Y(_06338_));
 sky130_fd_sc_hd__and2_1 _13775_ (.A(_06320_),
    .B(_06322_),
    .X(_06339_));
 sky130_fd_sc_hd__o21a_1 _13776_ (.A1(_06339_),
    .A2(_06326_),
    .B1(_06325_),
    .X(_06341_));
 sky130_fd_sc_hd__nor2_1 _13777_ (.A(_06339_),
    .B(_06327_),
    .Y(_06342_));
 sky130_fd_sc_hd__a211o_1 _13778_ (.A1(_06335_),
    .A2(_06338_),
    .B1(_06341_),
    .C1(_06342_),
    .X(_06343_));
 sky130_fd_sc_hd__nor2_1 _13779_ (.A(_06332_),
    .B(_06333_),
    .Y(_06344_));
 sky130_fd_sc_hd__nor2_1 _13780_ (.A(_06334_),
    .B(_06344_),
    .Y(_06345_));
 sky130_fd_sc_hd__o22a_1 _13781_ (.A1(_06334_),
    .A2(_06338_),
    .B1(_06345_),
    .B2(_06337_),
    .X(_06346_));
 sky130_fd_sc_hd__o21ai_1 _13782_ (.A1(_05884_),
    .A2(_05889_),
    .B1(_05885_),
    .Y(_06347_));
 sky130_fd_sc_hd__or2b_1 _13783_ (.A(_06346_),
    .B_N(_06347_),
    .X(_06348_));
 sky130_fd_sc_hd__or2_1 _13784_ (.A(_05891_),
    .B(_05894_),
    .X(_06349_));
 sky130_fd_sc_hd__xor2_1 _13785_ (.A(_06346_),
    .B(_06347_),
    .X(_06350_));
 sky130_fd_sc_hd__a21o_1 _13786_ (.A1(_06349_),
    .A2(_05897_),
    .B1(_06350_),
    .X(_06352_));
 sky130_fd_sc_hd__nand2_1 _13787_ (.A(_06348_),
    .B(_06352_),
    .Y(_06353_));
 sky130_fd_sc_hd__o211a_1 _13788_ (.A1(_06341_),
    .A2(_06342_),
    .B1(_06335_),
    .C1(_06338_),
    .X(_06354_));
 sky130_fd_sc_hd__a21o_1 _13789_ (.A1(_06343_),
    .A2(_06353_),
    .B1(_06354_),
    .X(_06355_));
 sky130_fd_sc_hd__and2_1 _13790_ (.A(_06331_),
    .B(_06355_),
    .X(_06356_));
 sky130_fd_sc_hd__nor2_1 _13791_ (.A(_06292_),
    .B(_06312_),
    .Y(_06357_));
 sky130_fd_sc_hd__nor2_1 _13792_ (.A(_06311_),
    .B(_06357_),
    .Y(_06358_));
 sky130_fd_sc_hd__o21a_1 _13793_ (.A1(_06328_),
    .A2(_06356_),
    .B1(_06358_),
    .X(_06359_));
 sky130_fd_sc_hd__nor3_1 _13794_ (.A(_06289_),
    .B(_06262_),
    .C(_06287_),
    .Y(_06360_));
 sky130_fd_sc_hd__nor2_1 _13795_ (.A(_06290_),
    .B(_06360_),
    .Y(_06361_));
 sky130_fd_sc_hd__o21a_1 _13796_ (.A1(_06311_),
    .A2(_06359_),
    .B1(_06361_),
    .X(_06363_));
 sky130_fd_sc_hd__nor4_1 _13797_ (.A(_06242_),
    .B(_06253_),
    .C(_06290_),
    .D(_06363_),
    .Y(_06364_));
 sky130_fd_sc_hd__and4_1 _13798_ (.A(_02188_),
    .B(_02190_),
    .C(_03684_),
    .D(_03680_),
    .X(_06365_));
 sky130_fd_sc_hd__and4_1 _13799_ (.A(_02187_),
    .B(_02189_),
    .C(_03686_),
    .D(_03683_),
    .X(_06366_));
 sky130_fd_sc_hd__nand2_1 _13800_ (.A(_02187_),
    .B(_03682_),
    .Y(_06367_));
 sky130_fd_sc_hd__a21boi_1 _13801_ (.A1(_02189_),
    .A2(_03686_),
    .B1_N(_06367_),
    .Y(_06368_));
 sky130_fd_sc_hd__nor2_1 _13802_ (.A(_06366_),
    .B(_06368_),
    .Y(_06369_));
 sky130_fd_sc_hd__and3_1 _13803_ (.A(_03414_),
    .B(_03679_),
    .C(_06369_),
    .X(_06370_));
 sky130_fd_sc_hd__a22oi_1 _13804_ (.A1(_02190_),
    .A2(_03684_),
    .B1(_03680_),
    .B2(_02188_),
    .Y(_06371_));
 sky130_fd_sc_hd__nor2_1 _13805_ (.A(_06365_),
    .B(_06371_),
    .Y(_06372_));
 sky130_fd_sc_hd__o21a_1 _13806_ (.A1(_06366_),
    .A2(_06370_),
    .B1(_06372_),
    .X(_06374_));
 sky130_fd_sc_hd__and3_1 _13807_ (.A(_02190_),
    .B(_03699_),
    .C(_06367_),
    .X(_06375_));
 sky130_fd_sc_hd__and2_1 _13808_ (.A(_06374_),
    .B(_06375_),
    .X(_06376_));
 sky130_fd_sc_hd__and4_1 _13809_ (.A(_02187_),
    .B(_02189_),
    .C(_01954_),
    .D(_03686_),
    .X(_06377_));
 sky130_fd_sc_hd__a22oi_1 _13810_ (.A1(_02189_),
    .A2(_01955_),
    .B1(_03686_),
    .B2(_02188_),
    .Y(_06378_));
 sky130_fd_sc_hd__and4bb_1 _13811_ (.A_N(_06377_),
    .B_N(_06378_),
    .C(_01400_),
    .D(_03683_),
    .X(_06379_));
 sky130_fd_sc_hd__nor2_1 _13812_ (.A(_06377_),
    .B(_06379_),
    .Y(_06380_));
 sky130_fd_sc_hd__a21oi_1 _13813_ (.A1(_03414_),
    .A2(_03679_),
    .B1(_06369_),
    .Y(_06381_));
 sky130_fd_sc_hd__or3_1 _13814_ (.A(_06370_),
    .B(_06380_),
    .C(_06381_),
    .X(_06382_));
 sky130_fd_sc_hd__nor3_1 _13815_ (.A(_06366_),
    .B(_06370_),
    .C(_06372_),
    .Y(_06383_));
 sky130_fd_sc_hd__nor2_1 _13816_ (.A(_06374_),
    .B(_06383_),
    .Y(_06385_));
 sky130_fd_sc_hd__and2b_1 _13817_ (.A_N(_06382_),
    .B(_06385_),
    .X(_06386_));
 sky130_fd_sc_hd__and3_1 _13818_ (.A(_01400_),
    .B(_02187_),
    .C(_03686_),
    .X(_06387_));
 sky130_fd_sc_hd__a22o_1 _13819_ (.A1(_02187_),
    .A2(_01955_),
    .B1(_03686_),
    .B2(_01400_),
    .X(_06388_));
 sky130_fd_sc_hd__a21bo_1 _13820_ (.A1(_01955_),
    .A2(_06387_),
    .B1_N(_06388_),
    .X(_06389_));
 sky130_fd_sc_hd__nand2_1 _13821_ (.A(_04714_),
    .B(_03683_),
    .Y(_06390_));
 sky130_fd_sc_hd__xnor2_1 _13822_ (.A(_06389_),
    .B(_06390_),
    .Y(_06391_));
 sky130_fd_sc_hd__nor2_1 _13823_ (.A(_05935_),
    .B(_06391_),
    .Y(_06392_));
 sky130_fd_sc_hd__o2bb2a_1 _13824_ (.A1_N(_03414_),
    .A2_N(_03683_),
    .B1(_06377_),
    .B2(_06378_),
    .X(_06393_));
 sky130_fd_sc_hd__or2_1 _13825_ (.A(_06379_),
    .B(_06393_),
    .X(_06394_));
 sky130_fd_sc_hd__a32o_1 _13826_ (.A1(_00460_),
    .A2(_03683_),
    .A3(_06388_),
    .B1(_06387_),
    .B2(_01955_),
    .X(_06396_));
 sky130_fd_sc_hd__and3_1 _13827_ (.A(_01066_),
    .B(_03679_),
    .C(_06396_),
    .X(_06397_));
 sky130_fd_sc_hd__a21oi_1 _13828_ (.A1(_04714_),
    .A2(_03680_),
    .B1(_06396_),
    .Y(_06398_));
 sky130_fd_sc_hd__nor2_1 _13829_ (.A(_06397_),
    .B(_06398_),
    .Y(_06399_));
 sky130_fd_sc_hd__xnor2_1 _13830_ (.A(_06394_),
    .B(_06399_),
    .Y(_06400_));
 sky130_fd_sc_hd__nand2_1 _13831_ (.A(_06392_),
    .B(_06400_),
    .Y(_06401_));
 sky130_fd_sc_hd__and2b_1 _13832_ (.A_N(_06394_),
    .B(_06399_),
    .X(_06402_));
 sky130_fd_sc_hd__o21ai_1 _13833_ (.A1(_06370_),
    .A2(_06381_),
    .B1(_06380_),
    .Y(_06403_));
 sky130_fd_sc_hd__and2_1 _13834_ (.A(_06382_),
    .B(_06403_),
    .X(_06404_));
 sky130_fd_sc_hd__o21ai_1 _13835_ (.A1(_06397_),
    .A2(_06402_),
    .B1(_06404_),
    .Y(_06405_));
 sky130_fd_sc_hd__or3_1 _13836_ (.A(_06397_),
    .B(_06402_),
    .C(_06404_),
    .X(_06407_));
 sky130_fd_sc_hd__nand2_1 _13837_ (.A(_06405_),
    .B(_06407_),
    .Y(_06408_));
 sky130_fd_sc_hd__o21a_1 _13838_ (.A1(_06401_),
    .A2(_06408_),
    .B1(_06405_),
    .X(_06409_));
 sky130_fd_sc_hd__xnor2_1 _13839_ (.A(_06382_),
    .B(_06385_),
    .Y(_06410_));
 sky130_fd_sc_hd__and2b_1 _13840_ (.A_N(_06409_),
    .B(_06410_),
    .X(_06411_));
 sky130_fd_sc_hd__nor2_1 _13841_ (.A(_06374_),
    .B(_06375_),
    .Y(_06412_));
 sky130_fd_sc_hd__nor2_1 _13842_ (.A(_06376_),
    .B(_06412_),
    .Y(_06413_));
 sky130_fd_sc_hd__o21a_1 _13843_ (.A1(_06386_),
    .A2(_06411_),
    .B1(_06413_),
    .X(_06414_));
 sky130_fd_sc_hd__and2b_1 _13844_ (.A_N(_06410_),
    .B(_06409_),
    .X(_06415_));
 sky130_fd_sc_hd__nor2_1 _13845_ (.A(_06411_),
    .B(_06415_),
    .Y(_06416_));
 sky130_fd_sc_hd__nor2_1 _13846_ (.A(_05902_),
    .B(_05905_),
    .Y(_06418_));
 sky130_fd_sc_hd__and3_1 _13847_ (.A(_02189_),
    .B(_03783_),
    .C(_05370_),
    .X(_06419_));
 sky130_fd_sc_hd__nand2_1 _13848_ (.A(_06418_),
    .B(_06419_),
    .Y(_06420_));
 sky130_fd_sc_hd__xor2_1 _13849_ (.A(_06418_),
    .B(_06419_),
    .X(_06421_));
 sky130_fd_sc_hd__o21ai_1 _13850_ (.A1(_05907_),
    .A2(_05911_),
    .B1(_06421_),
    .Y(_06422_));
 sky130_fd_sc_hd__and3_1 _13851_ (.A(_05904_),
    .B(_06420_),
    .C(_06422_),
    .X(_06423_));
 sky130_fd_sc_hd__nor2_1 _13852_ (.A(_05916_),
    .B(_05919_),
    .Y(_06424_));
 sky130_fd_sc_hd__and3_1 _13853_ (.A(_01517_),
    .B(_03679_),
    .C(_05386_),
    .X(_06425_));
 sky130_fd_sc_hd__nand2_1 _13854_ (.A(_06424_),
    .B(_06425_),
    .Y(_06426_));
 sky130_fd_sc_hd__xor2_1 _13855_ (.A(_06424_),
    .B(_06425_),
    .X(_06427_));
 sky130_fd_sc_hd__o21ai_1 _13856_ (.A1(_05921_),
    .A2(_05926_),
    .B1(_06427_),
    .Y(_06429_));
 sky130_fd_sc_hd__and3_1 _13857_ (.A(_05918_),
    .B(_06426_),
    .C(_06429_),
    .X(_06430_));
 sky130_fd_sc_hd__nor2_1 _13858_ (.A(_06423_),
    .B(_06430_),
    .Y(_06431_));
 sky130_fd_sc_hd__xor2_1 _13859_ (.A(_06401_),
    .B(_06408_),
    .X(_06432_));
 sky130_fd_sc_hd__and3_1 _13860_ (.A(_06416_),
    .B(_06431_),
    .C(_06432_),
    .X(_06433_));
 sky130_fd_sc_hd__and2_1 _13861_ (.A(_06431_),
    .B(_06432_),
    .X(_06434_));
 sky130_fd_sc_hd__nor2_1 _13862_ (.A(_06431_),
    .B(_06432_),
    .Y(_06435_));
 sky130_fd_sc_hd__nor2_1 _13863_ (.A(_06434_),
    .B(_06435_),
    .Y(_06436_));
 sky130_fd_sc_hd__or3_1 _13864_ (.A(_05907_),
    .B(_05911_),
    .C(_06421_),
    .X(_06437_));
 sky130_fd_sc_hd__and2_1 _13865_ (.A(_06422_),
    .B(_06437_),
    .X(_06438_));
 sky130_fd_sc_hd__or3_1 _13866_ (.A(_05921_),
    .B(_05926_),
    .C(_06427_),
    .X(_06440_));
 sky130_fd_sc_hd__and2_1 _13867_ (.A(_06429_),
    .B(_06440_),
    .X(_06441_));
 sky130_fd_sc_hd__nand2_1 _13868_ (.A(_06438_),
    .B(_06441_),
    .Y(_06442_));
 sky130_fd_sc_hd__and2_1 _13869_ (.A(_06423_),
    .B(_06430_),
    .X(_06443_));
 sky130_fd_sc_hd__or2_1 _13870_ (.A(_06431_),
    .B(_06443_),
    .X(_06444_));
 sky130_fd_sc_hd__nand2_1 _13871_ (.A(_06442_),
    .B(_06444_),
    .Y(_06445_));
 sky130_fd_sc_hd__or2_1 _13872_ (.A(_06392_),
    .B(_06400_),
    .X(_06446_));
 sky130_fd_sc_hd__and2_1 _13873_ (.A(_06401_),
    .B(_06446_),
    .X(_06447_));
 sky130_fd_sc_hd__nor2_1 _13874_ (.A(_06442_),
    .B(_06444_),
    .Y(_06448_));
 sky130_fd_sc_hd__or2_1 _13875_ (.A(_06447_),
    .B(_06448_),
    .X(_06449_));
 sky130_fd_sc_hd__and3_1 _13876_ (.A(_06436_),
    .B(_06445_),
    .C(_06449_),
    .X(_06451_));
 sky130_fd_sc_hd__a21oi_1 _13877_ (.A1(_06445_),
    .A2(_06449_),
    .B1(_06436_),
    .Y(_06452_));
 sky130_fd_sc_hd__nor2_1 _13878_ (.A(_06451_),
    .B(_06452_),
    .Y(_06453_));
 sky130_fd_sc_hd__nand2_1 _13879_ (.A(_05913_),
    .B(_05927_),
    .Y(_06454_));
 sky130_fd_sc_hd__xnor2_1 _13880_ (.A(_06438_),
    .B(_06441_),
    .Y(_06455_));
 sky130_fd_sc_hd__and2_1 _13881_ (.A(_06454_),
    .B(_06455_),
    .X(_06456_));
 sky130_fd_sc_hd__inv_2 _13882_ (.A(_06456_),
    .Y(_06457_));
 sky130_fd_sc_hd__and2_1 _13883_ (.A(_05935_),
    .B(_06391_),
    .X(_06458_));
 sky130_fd_sc_hd__or2_1 _13884_ (.A(_06392_),
    .B(_06458_),
    .X(_06459_));
 sky130_fd_sc_hd__o21ai_2 _13885_ (.A1(_06454_),
    .A2(_06455_),
    .B1(_06459_),
    .Y(_06460_));
 sky130_fd_sc_hd__and2_1 _13886_ (.A(_06442_),
    .B(_06444_),
    .X(_06462_));
 sky130_fd_sc_hd__o21a_1 _13887_ (.A1(_06462_),
    .A2(_06448_),
    .B1(_06447_),
    .X(_06463_));
 sky130_fd_sc_hd__nor2_1 _13888_ (.A(_06462_),
    .B(_06449_),
    .Y(_06464_));
 sky130_fd_sc_hd__a211o_1 _13889_ (.A1(_06457_),
    .A2(_06460_),
    .B1(_06463_),
    .C1(_06464_),
    .X(_06465_));
 sky130_fd_sc_hd__nor2_1 _13890_ (.A(_06454_),
    .B(_06455_),
    .Y(_06466_));
 sky130_fd_sc_hd__nor2_1 _13891_ (.A(_06456_),
    .B(_06466_),
    .Y(_06467_));
 sky130_fd_sc_hd__o22a_1 _13892_ (.A1(_06456_),
    .A2(_06460_),
    .B1(_06467_),
    .B2(_06459_),
    .X(_06468_));
 sky130_fd_sc_hd__a21bo_1 _13893_ (.A1(_05929_),
    .A2(_05936_),
    .B1_N(_05930_),
    .X(_06469_));
 sky130_fd_sc_hd__or2b_1 _13894_ (.A(_06468_),
    .B_N(_06469_),
    .X(_06470_));
 sky130_fd_sc_hd__or2_1 _13895_ (.A(_05937_),
    .B(_05940_),
    .X(_06471_));
 sky130_fd_sc_hd__or3_1 _13896_ (.A(_05363_),
    .B(_05405_),
    .C(_05941_),
    .X(_06473_));
 sky130_fd_sc_hd__xor2_1 _13897_ (.A(_06468_),
    .B(_06469_),
    .X(_06474_));
 sky130_fd_sc_hd__a21o_1 _13898_ (.A1(_06471_),
    .A2(_06473_),
    .B1(_06474_),
    .X(_06475_));
 sky130_fd_sc_hd__nand2_1 _13899_ (.A(_06470_),
    .B(_06475_),
    .Y(_06476_));
 sky130_fd_sc_hd__o211a_1 _13900_ (.A1(_06463_),
    .A2(_06464_),
    .B1(_06457_),
    .C1(_06460_),
    .X(_06477_));
 sky130_fd_sc_hd__a21o_1 _13901_ (.A1(_06465_),
    .A2(_06476_),
    .B1(_06477_),
    .X(_06478_));
 sky130_fd_sc_hd__and2_1 _13902_ (.A(_06453_),
    .B(_06478_),
    .X(_06479_));
 sky130_fd_sc_hd__nor2_1 _13903_ (.A(_06416_),
    .B(_06434_),
    .Y(_06480_));
 sky130_fd_sc_hd__nor2_1 _13904_ (.A(_06433_),
    .B(_06480_),
    .Y(_06481_));
 sky130_fd_sc_hd__o21a_1 _13905_ (.A1(_06451_),
    .A2(_06479_),
    .B1(_06481_),
    .X(_06482_));
 sky130_fd_sc_hd__nor3_1 _13906_ (.A(_06413_),
    .B(_06386_),
    .C(_06411_),
    .Y(_06484_));
 sky130_fd_sc_hd__nor2_1 _13907_ (.A(_06414_),
    .B(_06484_),
    .Y(_06485_));
 sky130_fd_sc_hd__o21a_1 _13908_ (.A1(_06433_),
    .A2(_06482_),
    .B1(_06485_),
    .X(_06486_));
 sky130_fd_sc_hd__nor4_1 _13909_ (.A(_06365_),
    .B(_06376_),
    .C(_06414_),
    .D(_06486_),
    .Y(_06487_));
 sky130_fd_sc_hd__nor2_1 _13910_ (.A(net137),
    .B(net136),
    .Y(_06488_));
 sky130_fd_sc_hd__or3_1 _13911_ (.A(_06234_),
    .B(_06201_),
    .C(_06231_),
    .X(_06489_));
 sky130_fd_sc_hd__and2_1 _13912_ (.A(_06235_),
    .B(_06489_),
    .X(_06490_));
 sky130_fd_sc_hd__and2_1 _13913_ (.A(_06488_),
    .B(_06490_),
    .X(_06491_));
 sky130_fd_sc_hd__mux2_2 _13914_ (.A0(_06240_),
    .A1(_06188_),
    .S(_06491_),
    .X(_06492_));
 sky130_fd_sc_hd__nor2_1 _13915_ (.A(_06488_),
    .B(_06490_),
    .Y(_06493_));
 sky130_fd_sc_hd__nor3_1 _13916_ (.A(_06361_),
    .B(_06311_),
    .C(_06359_),
    .Y(_06495_));
 sky130_fd_sc_hd__nor2_1 _13917_ (.A(_06363_),
    .B(_06495_),
    .Y(_06496_));
 sky130_fd_sc_hd__nor3_1 _13918_ (.A(_06485_),
    .B(_06433_),
    .C(_06482_),
    .Y(_06497_));
 sky130_fd_sc_hd__nor2_1 _13919_ (.A(_06486_),
    .B(_06497_),
    .Y(_06498_));
 sky130_fd_sc_hd__nand2_1 _13920_ (.A(_06496_),
    .B(_06498_),
    .Y(_06499_));
 sky130_fd_sc_hd__xnor2_1 _13921_ (.A(net137),
    .B(net136),
    .Y(_06500_));
 sky130_fd_sc_hd__and2_1 _13922_ (.A(_06499_),
    .B(_06500_),
    .X(_06501_));
 sky130_fd_sc_hd__xnor2_1 _13923_ (.A(_06203_),
    .B(_06229_),
    .Y(_06502_));
 sky130_fd_sc_hd__o21a_1 _13924_ (.A1(_06499_),
    .A2(_06500_),
    .B1(_06502_),
    .X(_06503_));
 sky130_fd_sc_hd__nor4_1 _13925_ (.A(_06491_),
    .B(_06493_),
    .C(_06501_),
    .D(_06503_),
    .Y(_06504_));
 sky130_fd_sc_hd__o22a_1 _13926_ (.A1(_06491_),
    .A2(_06493_),
    .B1(_06501_),
    .B2(_06503_),
    .X(_06506_));
 sky130_fd_sc_hd__or2_2 _13927_ (.A(net134),
    .B(_06506_),
    .X(_06507_));
 sky130_fd_sc_hd__nor2_2 _13928_ (.A(_06226_),
    .B(_06228_),
    .Y(_06508_));
 sky130_fd_sc_hd__xnor2_4 _13929_ (.A(_06220_),
    .B(_06508_),
    .Y(_06509_));
 sky130_fd_sc_hd__nor3_1 _13930_ (.A(_06358_),
    .B(_06328_),
    .C(_06356_),
    .Y(_06510_));
 sky130_fd_sc_hd__nor2_1 _13931_ (.A(_06359_),
    .B(_06510_),
    .Y(_06511_));
 sky130_fd_sc_hd__nor3_1 _13932_ (.A(_06481_),
    .B(_06451_),
    .C(_06479_),
    .Y(_06512_));
 sky130_fd_sc_hd__nor2_1 _13933_ (.A(_06482_),
    .B(_06512_),
    .Y(_06513_));
 sky130_fd_sc_hd__nand2_1 _13934_ (.A(_06511_),
    .B(_06513_),
    .Y(_06514_));
 sky130_fd_sc_hd__or2_1 _13935_ (.A(_06496_),
    .B(_06498_),
    .X(_06515_));
 sky130_fd_sc_hd__nand2_1 _13936_ (.A(_06499_),
    .B(_06515_),
    .Y(_06517_));
 sky130_fd_sc_hd__nor2_1 _13937_ (.A(_06514_),
    .B(_06517_),
    .Y(_06518_));
 sky130_fd_sc_hd__nand2_1 _13938_ (.A(_06514_),
    .B(_06517_),
    .Y(_06519_));
 sky130_fd_sc_hd__and2b_1 _13939_ (.A_N(_06518_),
    .B(_06519_),
    .X(_06520_));
 sky130_fd_sc_hd__xnor2_4 _13940_ (.A(_06509_),
    .B(_06520_),
    .Y(_06521_));
 sky130_fd_sc_hd__and2_1 _13941_ (.A(_06226_),
    .B(_06228_),
    .X(_06522_));
 sky130_fd_sc_hd__nor2_1 _13942_ (.A(_06508_),
    .B(_06522_),
    .Y(_06523_));
 sky130_fd_sc_hd__xor2_2 _13943_ (.A(_06331_),
    .B(_06355_),
    .X(_06524_));
 sky130_fd_sc_hd__xor2_2 _13944_ (.A(_06453_),
    .B(_06478_),
    .X(_06525_));
 sky130_fd_sc_hd__nand2_1 _13945_ (.A(_06524_),
    .B(_06525_),
    .Y(_06526_));
 sky130_fd_sc_hd__or2_1 _13946_ (.A(_06511_),
    .B(_06513_),
    .X(_06528_));
 sky130_fd_sc_hd__nand2_1 _13947_ (.A(_06514_),
    .B(_06528_),
    .Y(_06529_));
 sky130_fd_sc_hd__nor2_1 _13948_ (.A(_06526_),
    .B(_06529_),
    .Y(_06530_));
 sky130_fd_sc_hd__and2_1 _13949_ (.A(_06526_),
    .B(_06529_),
    .X(_06531_));
 sky130_fd_sc_hd__o21ba_2 _13950_ (.A1(_06523_),
    .A2(_06530_),
    .B1_N(_06531_),
    .X(_06532_));
 sky130_fd_sc_hd__xnor2_4 _13951_ (.A(_06521_),
    .B(_06532_),
    .Y(_06533_));
 sky130_fd_sc_hd__and2b_1 _13952_ (.A_N(_06225_),
    .B(_06224_),
    .X(_06534_));
 sky130_fd_sc_hd__xnor2_1 _13953_ (.A(_06221_),
    .B(_06534_),
    .Y(_06535_));
 sky130_fd_sc_hd__and2b_1 _13954_ (.A_N(_06354_),
    .B(_06343_),
    .X(_06536_));
 sky130_fd_sc_hd__xnor2_1 _13955_ (.A(_06353_),
    .B(_06536_),
    .Y(_06537_));
 sky130_fd_sc_hd__and2b_1 _13956_ (.A_N(_06477_),
    .B(_06465_),
    .X(_06539_));
 sky130_fd_sc_hd__xnor2_2 _13957_ (.A(_06476_),
    .B(_06539_),
    .Y(_06540_));
 sky130_fd_sc_hd__or2_1 _13958_ (.A(_06537_),
    .B(_06540_),
    .X(_06541_));
 sky130_fd_sc_hd__xnor2_1 _13959_ (.A(_06524_),
    .B(_06525_),
    .Y(_06542_));
 sky130_fd_sc_hd__nand2_1 _13960_ (.A(_06541_),
    .B(_06542_),
    .Y(_06543_));
 sky130_fd_sc_hd__inv_2 _13961_ (.A(_06543_),
    .Y(_06544_));
 sky130_fd_sc_hd__nor2_1 _13962_ (.A(_06541_),
    .B(_06542_),
    .Y(_06545_));
 sky130_fd_sc_hd__nor2_1 _13963_ (.A(_06544_),
    .B(_06545_),
    .Y(_06546_));
 sky130_fd_sc_hd__xnor2_1 _13964_ (.A(_06535_),
    .B(_06546_),
    .Y(_06547_));
 sky130_fd_sc_hd__nand3_1 _13965_ (.A(_06349_),
    .B(_05897_),
    .C(_06350_),
    .Y(_06548_));
 sky130_fd_sc_hd__nand2_1 _13966_ (.A(_06352_),
    .B(_06548_),
    .Y(_06550_));
 sky130_fd_sc_hd__nand3_1 _13967_ (.A(_06471_),
    .B(_06473_),
    .C(_06474_),
    .Y(_06551_));
 sky130_fd_sc_hd__nand2_1 _13968_ (.A(_06475_),
    .B(_06551_),
    .Y(_06552_));
 sky130_fd_sc_hd__nor2_1 _13969_ (.A(_06550_),
    .B(_06552_),
    .Y(_06553_));
 sky130_fd_sc_hd__nand2_1 _13970_ (.A(_06537_),
    .B(_06540_),
    .Y(_06554_));
 sky130_fd_sc_hd__and2_1 _13971_ (.A(_06541_),
    .B(_06554_),
    .X(_06555_));
 sky130_fd_sc_hd__nor2_1 _13972_ (.A(_06553_),
    .B(_06555_),
    .Y(_06556_));
 sky130_fd_sc_hd__or2_1 _13973_ (.A(_06157_),
    .B(_06159_),
    .X(_06557_));
 sky130_fd_sc_hd__nand2_1 _13974_ (.A(_06160_),
    .B(_06557_),
    .Y(_06558_));
 sky130_fd_sc_hd__nand2_1 _13975_ (.A(_06553_),
    .B(_06555_),
    .Y(_06559_));
 sky130_fd_sc_hd__and2_1 _13976_ (.A(_06558_),
    .B(_06559_),
    .X(_06561_));
 sky130_fd_sc_hd__nor3_1 _13977_ (.A(_06547_),
    .B(_06556_),
    .C(_06561_),
    .Y(_06562_));
 sky130_fd_sc_hd__and2b_1 _13978_ (.A_N(_05947_),
    .B(_05952_),
    .X(_06563_));
 sky130_fd_sc_hd__and2_1 _13979_ (.A(_05951_),
    .B(_06156_),
    .X(_06564_));
 sky130_fd_sc_hd__or2_1 _13980_ (.A(_06157_),
    .B(_06564_),
    .X(_06565_));
 sky130_fd_sc_hd__and2_1 _13981_ (.A(_06550_),
    .B(_06552_),
    .X(_06566_));
 sky130_fd_sc_hd__nor2_1 _13982_ (.A(_06553_),
    .B(_06566_),
    .Y(_06567_));
 sky130_fd_sc_hd__and3_1 _13983_ (.A(_05898_),
    .B(_05942_),
    .C(_06567_),
    .X(_06568_));
 sky130_fd_sc_hd__a21oi_1 _13984_ (.A1(_05898_),
    .A2(_05942_),
    .B1(_06567_),
    .Y(_06569_));
 sky130_fd_sc_hd__nor2_1 _13985_ (.A(_06568_),
    .B(_06569_),
    .Y(_06570_));
 sky130_fd_sc_hd__xnor2_1 _13986_ (.A(_06565_),
    .B(_06570_),
    .Y(_06572_));
 sky130_fd_sc_hd__o21a_1 _13987_ (.A1(_05946_),
    .A2(_06563_),
    .B1(_06572_),
    .X(_06573_));
 sky130_fd_sc_hd__nor2_1 _13988_ (.A(_06565_),
    .B(_06569_),
    .Y(_06574_));
 sky130_fd_sc_hd__and2b_1 _13989_ (.A_N(_06556_),
    .B(_06559_),
    .X(_06575_));
 sky130_fd_sc_hd__xnor2_1 _13990_ (.A(_06558_),
    .B(_06575_),
    .Y(_06576_));
 sky130_fd_sc_hd__o21ai_2 _13991_ (.A1(_06568_),
    .A2(_06574_),
    .B1(_06576_),
    .Y(_06577_));
 sky130_fd_sc_hd__inv_2 _13992_ (.A(_06577_),
    .Y(_06578_));
 sky130_fd_sc_hd__nor3_1 _13993_ (.A(_05946_),
    .B(_06563_),
    .C(_06572_),
    .Y(_06579_));
 sky130_fd_sc_hd__nor2_1 _13994_ (.A(_06573_),
    .B(_06579_),
    .Y(_06580_));
 sky130_fd_sc_hd__o211a_1 _13995_ (.A1(_05417_),
    .A2(_05954_),
    .B1(_05955_),
    .C1(_06580_),
    .X(_06581_));
 sky130_fd_sc_hd__nor3_1 _13996_ (.A(_06576_),
    .B(_06568_),
    .C(_06574_),
    .Y(_06583_));
 sky130_fd_sc_hd__inv_2 _13997_ (.A(_06583_),
    .Y(_06584_));
 sky130_fd_sc_hd__o21a_1 _13998_ (.A1(_06556_),
    .A2(_06561_),
    .B1(_06547_),
    .X(_06585_));
 sky130_fd_sc_hd__nor2_1 _13999_ (.A(_06562_),
    .B(_06585_),
    .Y(_06586_));
 sky130_fd_sc_hd__o311a_1 _14000_ (.A1(_06573_),
    .A2(_06578_),
    .A3(_06581_),
    .B1(_06584_),
    .C1(_06586_),
    .X(_06587_));
 sky130_fd_sc_hd__o21ai_1 _14001_ (.A1(_06531_),
    .A2(_06530_),
    .B1(_06523_),
    .Y(_06588_));
 sky130_fd_sc_hd__or3_1 _14002_ (.A(_06531_),
    .B(_06523_),
    .C(_06530_),
    .X(_06589_));
 sky130_fd_sc_hd__and2_1 _14003_ (.A(_06588_),
    .B(_06589_),
    .X(_06590_));
 sky130_fd_sc_hd__o21ai_1 _14004_ (.A1(_06535_),
    .A2(_06545_),
    .B1(_06543_),
    .Y(_06591_));
 sky130_fd_sc_hd__nor2_1 _14005_ (.A(_06590_),
    .B(_06591_),
    .Y(_06592_));
 sky130_fd_sc_hd__and3_1 _14006_ (.A(_06588_),
    .B(_06589_),
    .C(_06591_),
    .X(_06594_));
 sky130_fd_sc_hd__inv_2 _14007_ (.A(_06594_),
    .Y(_06595_));
 sky130_fd_sc_hd__o31a_2 _14008_ (.A1(net132),
    .A2(_06587_),
    .A3(_06592_),
    .B1(_06595_),
    .X(_06596_));
 sky130_fd_sc_hd__and2b_1 _14009_ (.A_N(_06521_),
    .B(_06532_),
    .X(_06597_));
 sky130_fd_sc_hd__a21oi_4 _14010_ (.A1(_06533_),
    .A2(_06596_),
    .B1(_06597_),
    .Y(_06598_));
 sky130_fd_sc_hd__a21oi_1 _14011_ (.A1(_06509_),
    .A2(_06519_),
    .B1(_06518_),
    .Y(_06599_));
 sky130_fd_sc_hd__nor2_1 _14012_ (.A(_06499_),
    .B(_06500_),
    .Y(_06600_));
 sky130_fd_sc_hd__nor2_1 _14013_ (.A(_06501_),
    .B(_06600_),
    .Y(_06601_));
 sky130_fd_sc_hd__xnor2_1 _14014_ (.A(_06502_),
    .B(_06601_),
    .Y(_06602_));
 sky130_fd_sc_hd__xnor2_1 _14015_ (.A(_06599_),
    .B(_06602_),
    .Y(_06603_));
 sky130_fd_sc_hd__inv_2 _14016_ (.A(_06603_),
    .Y(_06605_));
 sky130_fd_sc_hd__or2b_1 _14017_ (.A(_06599_),
    .B_N(_06602_),
    .X(_06606_));
 sky130_fd_sc_hd__o21a_4 _14018_ (.A1(_06598_),
    .A2(_06605_),
    .B1(_06606_),
    .X(_06607_));
 sky130_fd_sc_hd__nor2_1 _14019_ (.A(_06491_),
    .B(_06504_),
    .Y(_06608_));
 sky130_fd_sc_hd__o32a_2 _14020_ (.A1(_06492_),
    .A2(_06507_),
    .A3(_06607_),
    .B1(_06608_),
    .B2(_06240_),
    .X(_06609_));
 sky130_fd_sc_hd__xnor2_4 _14021_ (.A(_06238_),
    .B(_06609_),
    .Y(_06610_));
 sky130_fd_sc_hd__nor2_1 _14022_ (.A(_05424_),
    .B(_05960_),
    .Y(_06611_));
 sky130_fd_sc_hd__o21a_1 _14023_ (.A1(_05851_),
    .A2(_05421_),
    .B1(_05958_),
    .X(_06612_));
 sky130_fd_sc_hd__a21o_1 _14024_ (.A1(_05750_),
    .A2(_06611_),
    .B1(_06612_),
    .X(_06613_));
 sky130_fd_sc_hd__a31o_1 _14025_ (.A1(_05810_),
    .A2(_05811_),
    .A3(_05812_),
    .B1(_05835_),
    .X(_06614_));
 sky130_fd_sc_hd__nand2_1 _14026_ (.A(_05648_),
    .B(_06611_),
    .Y(_06616_));
 sky130_fd_sc_hd__a21oi_2 _14027_ (.A1(_05839_),
    .A2(_06614_),
    .B1(_06616_),
    .Y(_06617_));
 sky130_fd_sc_hd__o21ai_2 _14028_ (.A1(_05417_),
    .A2(_05954_),
    .B1(_05955_),
    .Y(_06618_));
 sky130_fd_sc_hd__xor2_2 _14029_ (.A(_06618_),
    .B(_06580_),
    .X(_06619_));
 sky130_fd_sc_hd__inv_2 _14030_ (.A(_06619_),
    .Y(_06620_));
 sky130_fd_sc_hd__xnor2_4 _14031_ (.A(_06598_),
    .B(_06605_),
    .Y(_06621_));
 sky130_fd_sc_hd__xnor2_4 _14032_ (.A(_06507_),
    .B(_06607_),
    .Y(_06622_));
 sky130_fd_sc_hd__or2_1 _14033_ (.A(_06621_),
    .B(_06622_),
    .X(_06623_));
 sky130_fd_sc_hd__inv_2 _14034_ (.A(net133),
    .Y(_06624_));
 sky130_fd_sc_hd__a21o_1 _14035_ (.A1(_06624_),
    .A2(_06607_),
    .B1(_06506_),
    .X(_06625_));
 sky130_fd_sc_hd__xor2_4 _14036_ (.A(_06492_),
    .B(_06625_),
    .X(_06627_));
 sky130_fd_sc_hd__or2b_1 _14037_ (.A(_06623_),
    .B_N(_06627_),
    .X(_06628_));
 sky130_fd_sc_hd__o21ba_1 _14038_ (.A1(_06579_),
    .A2(_06618_),
    .B1_N(_06573_),
    .X(_06629_));
 sky130_fd_sc_hd__or3_2 _14039_ (.A(net135),
    .B(_06629_),
    .C(_06578_),
    .X(_06630_));
 sky130_fd_sc_hd__o21ai_1 _14040_ (.A1(net135),
    .A2(_06578_),
    .B1(_06629_),
    .Y(_06631_));
 sky130_fd_sc_hd__nand2_4 _14041_ (.A(_06630_),
    .B(_06631_),
    .Y(_06632_));
 sky130_fd_sc_hd__a21oi_1 _14042_ (.A1(_06629_),
    .A2(_06577_),
    .B1(net135),
    .Y(_06633_));
 sky130_fd_sc_hd__nor2_1 _14043_ (.A(_06586_),
    .B(_06633_),
    .Y(_06634_));
 sky130_fd_sc_hd__or2_2 _14044_ (.A(_06587_),
    .B(_06634_),
    .X(_06635_));
 sky130_fd_sc_hd__xnor2_2 _14045_ (.A(_06533_),
    .B(_06596_),
    .Y(_06636_));
 sky130_fd_sc_hd__nor2_1 _14046_ (.A(_06594_),
    .B(_06592_),
    .Y(_06638_));
 sky130_fd_sc_hd__inv_2 _14047_ (.A(net132),
    .Y(_06639_));
 sky130_fd_sc_hd__a31o_1 _14048_ (.A1(_06639_),
    .A2(_06577_),
    .A3(_06630_),
    .B1(_06585_),
    .X(_06640_));
 sky130_fd_sc_hd__xnor2_2 _14049_ (.A(_06638_),
    .B(_06640_),
    .Y(_06641_));
 sky130_fd_sc_hd__inv_2 _14050_ (.A(_06641_),
    .Y(_06642_));
 sky130_fd_sc_hd__or2_2 _14051_ (.A(_06636_),
    .B(_06642_),
    .X(_06643_));
 sky130_fd_sc_hd__or2_1 _14052_ (.A(_06635_),
    .B(_06643_),
    .X(_06644_));
 sky130_fd_sc_hd__or2_2 _14053_ (.A(_06632_),
    .B(_06644_),
    .X(_06645_));
 sky130_fd_sc_hd__nor2_1 _14054_ (.A(_06628_),
    .B(_06645_),
    .Y(_06646_));
 sky130_fd_sc_hd__o211a_1 _14055_ (.A1(_06613_),
    .A2(_06617_),
    .B1(_06620_),
    .C1(_06646_),
    .X(_06647_));
 sky130_fd_sc_hd__xnor2_4 _14056_ (.A(_06610_),
    .B(_06647_),
    .Y(net118));
 sky130_fd_sc_hd__or2_2 _14057_ (.A(_06238_),
    .B(_06609_),
    .X(_06649_));
 sky130_fd_sc_hd__inv_2 _14058_ (.A(_06111_),
    .Y(_06650_));
 sky130_fd_sc_hd__a21bo_1 _14059_ (.A1(_06062_),
    .A2(_06093_),
    .B1_N(_06061_),
    .X(_06651_));
 sky130_fd_sc_hd__and4_1 _14060_ (.A(_05969_),
    .B(_05985_),
    .C(_02743_),
    .D(_02742_),
    .X(_06652_));
 sky130_fd_sc_hd__a211o_1 _14061_ (.A1(_06085_),
    .A2(_06086_),
    .B1(_06090_),
    .C1(_06652_),
    .X(_06653_));
 sky130_fd_sc_hd__o21a_1 _14062_ (.A1(_06096_),
    .A2(_06651_),
    .B1(_06653_),
    .X(_06654_));
 sky130_fd_sc_hd__nor3_1 _14063_ (.A(_06096_),
    .B(_06653_),
    .C(_06651_),
    .Y(_06655_));
 sky130_fd_sc_hd__or2_1 _14064_ (.A(_06654_),
    .B(_06655_),
    .X(_06656_));
 sky130_fd_sc_hd__nand2_1 _14065_ (.A(_06099_),
    .B(_06656_),
    .Y(_06657_));
 sky130_fd_sc_hd__or2_1 _14066_ (.A(_06099_),
    .B(_06656_),
    .X(_06659_));
 sky130_fd_sc_hd__nand2_1 _14067_ (.A(_06657_),
    .B(_06659_),
    .Y(_06660_));
 sky130_fd_sc_hd__and2b_1 _14068_ (.A_N(_06108_),
    .B(_06079_),
    .X(_06661_));
 sky130_fd_sc_hd__a22oi_1 _14069_ (.A1(_06078_),
    .A2(_02743_),
    .B1(_02742_),
    .B2(_06075_),
    .Y(_06662_));
 sky130_fd_sc_hd__and4_1 _14070_ (.A(_06075_),
    .B(_06078_),
    .C(_02743_),
    .D(_02742_),
    .X(_06663_));
 sky130_fd_sc_hd__o2bb2a_1 _14071_ (.A1_N(_06077_),
    .A2_N(_04014_),
    .B1(_06662_),
    .B2(_06663_),
    .X(_06664_));
 sky130_fd_sc_hd__and4bb_1 _14072_ (.A_N(_06662_),
    .B_N(_06663_),
    .C(_06077_),
    .D(_04014_),
    .X(_06665_));
 sky130_fd_sc_hd__or2_1 _14073_ (.A(_06664_),
    .B(_06665_),
    .X(_06666_));
 sky130_fd_sc_hd__a41o_1 _14074_ (.A1(_06075_),
    .A2(_06077_),
    .A3(_06078_),
    .A4(_02743_),
    .B1(_06107_),
    .X(_06667_));
 sky130_fd_sc_hd__and3_1 _14075_ (.A(_06074_),
    .B(_04013_),
    .C(_06667_),
    .X(_06668_));
 sky130_fd_sc_hd__a21oi_1 _14076_ (.A1(_06074_),
    .A2(_04013_),
    .B1(_06667_),
    .Y(_06670_));
 sky130_fd_sc_hd__nor2_1 _14077_ (.A(_06668_),
    .B(_06670_),
    .Y(_06671_));
 sky130_fd_sc_hd__xnor2_1 _14078_ (.A(_06666_),
    .B(_06671_),
    .Y(_06672_));
 sky130_fd_sc_hd__nand2_1 _14079_ (.A(_06661_),
    .B(_06672_),
    .Y(_06673_));
 sky130_fd_sc_hd__or2_1 _14080_ (.A(_06661_),
    .B(_06672_),
    .X(_06674_));
 sky130_fd_sc_hd__nand2_1 _14081_ (.A(_06673_),
    .B(_06674_),
    .Y(_06675_));
 sky130_fd_sc_hd__xnor2_1 _14082_ (.A(_06660_),
    .B(_06675_),
    .Y(_06676_));
 sky130_fd_sc_hd__o21ai_1 _14083_ (.A1(_06102_),
    .A2(_06650_),
    .B1(_06676_),
    .Y(_06677_));
 sky130_fd_sc_hd__inv_2 _14084_ (.A(_06677_),
    .Y(_06678_));
 sky130_fd_sc_hd__nor3_1 _14085_ (.A(_06102_),
    .B(_06650_),
    .C(_06676_),
    .Y(_06679_));
 sky130_fd_sc_hd__nor2_2 _14086_ (.A(_06678_),
    .B(_06679_),
    .Y(_06681_));
 sky130_fd_sc_hd__a21o_2 _14087_ (.A1(_06116_),
    .A2(_06237_),
    .B1(_06115_),
    .X(_06682_));
 sky130_fd_sc_hd__xnor2_4 _14088_ (.A(_06681_),
    .B(_06682_),
    .Y(_06683_));
 sky130_fd_sc_hd__xnor2_4 _14089_ (.A(_06649_),
    .B(_06683_),
    .Y(_06684_));
 sky130_fd_sc_hd__nor2_1 _14090_ (.A(_05960_),
    .B(_06619_),
    .Y(_06685_));
 sky130_fd_sc_hd__nand2_1 _14091_ (.A(_05961_),
    .B(_06685_),
    .Y(_06686_));
 sky130_fd_sc_hd__o2bb2a_1 _14092_ (.A1_N(_05964_),
    .A2_N(_06685_),
    .B1(_06619_),
    .B2(_05959_),
    .X(_06687_));
 sky130_fd_sc_hd__or2b_1 _14093_ (.A(_06686_),
    .B_N(_05848_),
    .X(_06688_));
 sky130_fd_sc_hd__o311a_4 _14094_ (.A1(_05821_),
    .A2(_05842_),
    .A3(_06686_),
    .B1(_06687_),
    .C1(_06688_),
    .X(_06689_));
 sky130_fd_sc_hd__or2_1 _14095_ (.A(_06610_),
    .B(_06628_),
    .X(_06690_));
 sky130_fd_sc_hd__or3_4 _14096_ (.A(_06645_),
    .B(_06689_),
    .C(_06690_),
    .X(_06692_));
 sky130_fd_sc_hd__xor2_4 _14097_ (.A(_06684_),
    .B(_06692_),
    .X(net119));
 sky130_fd_sc_hd__nor2_1 _14098_ (.A(_06619_),
    .B(_06632_),
    .Y(_06693_));
 sky130_fd_sc_hd__and2_1 _14099_ (.A(_06611_),
    .B(_06693_),
    .X(_06694_));
 sky130_fd_sc_hd__and3_1 _14100_ (.A(_05648_),
    .B(_05679_),
    .C(_06694_),
    .X(_06695_));
 sky130_fd_sc_hd__a22o_1 _14101_ (.A1(_06612_),
    .A2(_06693_),
    .B1(_06694_),
    .B2(_05751_),
    .X(_06696_));
 sky130_fd_sc_hd__a21oi_4 _14102_ (.A1(_05825_),
    .A2(_06695_),
    .B1(_06696_),
    .Y(_06697_));
 sky130_fd_sc_hd__or2_1 _14103_ (.A(_06684_),
    .B(_06690_),
    .X(_06698_));
 sky130_fd_sc_hd__or3_4 _14104_ (.A(_06644_),
    .B(_06697_),
    .C(_06698_),
    .X(_06699_));
 sky130_fd_sc_hd__o21ba_1 _14105_ (.A1(_06666_),
    .A2(_06670_),
    .B1_N(_06668_),
    .X(_06700_));
 sky130_fd_sc_hd__nand2_1 _14106_ (.A(_02743_),
    .B(_04014_),
    .Y(_06702_));
 sky130_fd_sc_hd__a21boi_1 _14107_ (.A1(_06078_),
    .A2(_02742_),
    .B1_N(_06702_),
    .Y(_06703_));
 sky130_fd_sc_hd__and4_1 _14108_ (.A(_06078_),
    .B(_02743_),
    .C(_04014_),
    .D(_02742_),
    .X(_06704_));
 sky130_fd_sc_hd__nor2_1 _14109_ (.A(_06703_),
    .B(_06704_),
    .Y(_06705_));
 sky130_fd_sc_hd__nand2_1 _14110_ (.A(_06077_),
    .B(_04013_),
    .Y(_06706_));
 sky130_fd_sc_hd__xnor2_1 _14111_ (.A(_06705_),
    .B(_06706_),
    .Y(_06707_));
 sky130_fd_sc_hd__o21ai_1 _14112_ (.A1(_06663_),
    .A2(_06665_),
    .B1(_06707_),
    .Y(_06708_));
 sky130_fd_sc_hd__or3_1 _14113_ (.A(_06663_),
    .B(_06665_),
    .C(_06707_),
    .X(_06709_));
 sky130_fd_sc_hd__and2_1 _14114_ (.A(_06708_),
    .B(_06709_),
    .X(_06710_));
 sky130_fd_sc_hd__xnor2_1 _14115_ (.A(_06700_),
    .B(_06710_),
    .Y(_06711_));
 sky130_fd_sc_hd__xnor2_1 _14116_ (.A(_06673_),
    .B(_06711_),
    .Y(_06713_));
 sky130_fd_sc_hd__and2_1 _14117_ (.A(_06654_),
    .B(_06713_),
    .X(_06714_));
 sky130_fd_sc_hd__nor2_1 _14118_ (.A(_06654_),
    .B(_06713_),
    .Y(_06715_));
 sky130_fd_sc_hd__nor2_1 _14119_ (.A(_06714_),
    .B(_06715_),
    .Y(_06716_));
 sky130_fd_sc_hd__o21ai_1 _14120_ (.A1(_06099_),
    .A2(_06656_),
    .B1(_06675_),
    .Y(_06717_));
 sky130_fd_sc_hd__nand2_1 _14121_ (.A(_06657_),
    .B(_06717_),
    .Y(_06718_));
 sky130_fd_sc_hd__xnor2_1 _14122_ (.A(_06716_),
    .B(_06718_),
    .Y(_06719_));
 sky130_fd_sc_hd__inv_2 _14123_ (.A(_06719_),
    .Y(_06720_));
 sky130_fd_sc_hd__o21ai_1 _14124_ (.A1(_06679_),
    .A2(_06682_),
    .B1(_06677_),
    .Y(_06721_));
 sky130_fd_sc_hd__nor2_1 _14125_ (.A(_06720_),
    .B(_06721_),
    .Y(_06722_));
 sky130_fd_sc_hd__and2_1 _14126_ (.A(_06720_),
    .B(_06721_),
    .X(_06724_));
 sky130_fd_sc_hd__nor2_1 _14127_ (.A(_06722_),
    .B(_06724_),
    .Y(_06725_));
 sky130_fd_sc_hd__or3b_2 _14128_ (.A(_06649_),
    .B(_06683_),
    .C_N(_06725_),
    .X(_06726_));
 sky130_fd_sc_hd__o21bai_1 _14129_ (.A1(_06649_),
    .A2(_06683_),
    .B1_N(_06725_),
    .Y(_06727_));
 sky130_fd_sc_hd__nand2_2 _14130_ (.A(_06726_),
    .B(_06727_),
    .Y(_06728_));
 sky130_fd_sc_hd__xor2_4 _14131_ (.A(_06699_),
    .B(_06728_),
    .X(net121));
 sky130_fd_sc_hd__a31o_1 _14132_ (.A1(_06657_),
    .A2(_06717_),
    .A3(_06716_),
    .B1(_06722_),
    .X(_06729_));
 sky130_fd_sc_hd__a31o_1 _14133_ (.A1(_06077_),
    .A2(_04013_),
    .A3(_06705_),
    .B1(_06704_),
    .X(_06730_));
 sky130_fd_sc_hd__a22o_1 _14134_ (.A1(_04014_),
    .A2(_02742_),
    .B1(_04013_),
    .B2(_02743_),
    .X(_06731_));
 sky130_fd_sc_hd__nand4_1 _14135_ (.A(_02743_),
    .B(_04014_),
    .C(_02742_),
    .D(_04013_),
    .Y(_06732_));
 sky130_fd_sc_hd__nand2_1 _14136_ (.A(_06731_),
    .B(_06732_),
    .Y(_06734_));
 sky130_fd_sc_hd__xnor2_1 _14137_ (.A(_06730_),
    .B(_06734_),
    .Y(_06735_));
 sky130_fd_sc_hd__xnor2_1 _14138_ (.A(_06708_),
    .B(_06735_),
    .Y(_06736_));
 sky130_fd_sc_hd__and2b_1 _14139_ (.A_N(_06710_),
    .B(_06700_),
    .X(_06737_));
 sky130_fd_sc_hd__or2b_1 _14140_ (.A(_06700_),
    .B_N(_06710_),
    .X(_06738_));
 sky130_fd_sc_hd__o21a_1 _14141_ (.A1(_06673_),
    .A2(_06737_),
    .B1(_06738_),
    .X(_06739_));
 sky130_fd_sc_hd__and2b_1 _14142_ (.A_N(_06736_),
    .B(_06739_),
    .X(_06740_));
 sky130_fd_sc_hd__and2b_1 _14143_ (.A_N(_06739_),
    .B(_06736_),
    .X(_06741_));
 sky130_fd_sc_hd__nor2_1 _14144_ (.A(_06740_),
    .B(_06741_),
    .Y(_06742_));
 sky130_fd_sc_hd__nand2_1 _14145_ (.A(_06714_),
    .B(_06742_),
    .Y(_06743_));
 sky130_fd_sc_hd__or2_1 _14146_ (.A(_06714_),
    .B(_06742_),
    .X(_06745_));
 sky130_fd_sc_hd__nand2_1 _14147_ (.A(_06743_),
    .B(_06745_),
    .Y(_06746_));
 sky130_fd_sc_hd__or2b_1 _14148_ (.A(_06729_),
    .B_N(_06746_),
    .X(_06747_));
 sky130_fd_sc_hd__or2b_1 _14149_ (.A(_06746_),
    .B_N(_06729_),
    .X(_06748_));
 sky130_fd_sc_hd__nand2_1 _14150_ (.A(_06747_),
    .B(_06748_),
    .Y(_06749_));
 sky130_fd_sc_hd__or2_1 _14151_ (.A(_06726_),
    .B(_06749_),
    .X(_06750_));
 sky130_fd_sc_hd__nand2_1 _14152_ (.A(_06726_),
    .B(_06749_),
    .Y(_06751_));
 sky130_fd_sc_hd__nand2_2 _14153_ (.A(_06750_),
    .B(_06751_),
    .Y(_06752_));
 sky130_fd_sc_hd__or3_2 _14154_ (.A(_06619_),
    .B(_06632_),
    .C(_06635_),
    .X(_06753_));
 sky130_fd_sc_hd__nor2_1 _14155_ (.A(_05960_),
    .B(_06753_),
    .Y(_06754_));
 sky130_fd_sc_hd__o211ai_2 _14156_ (.A1(_05830_),
    .A2(_05833_),
    .B1(_05962_),
    .C1(_06754_),
    .Y(_06756_));
 sky130_fd_sc_hd__or2_1 _14157_ (.A(_05959_),
    .B(_06753_),
    .X(_06757_));
 sky130_fd_sc_hd__nand2_1 _14158_ (.A(_05965_),
    .B(_06754_),
    .Y(_06758_));
 sky130_fd_sc_hd__or2_2 _14159_ (.A(_06698_),
    .B(_06728_),
    .X(_06759_));
 sky130_fd_sc_hd__a311oi_4 _14160_ (.A1(_06756_),
    .A2(_06757_),
    .A3(_06758_),
    .B1(_06759_),
    .C1(_06643_),
    .Y(_06760_));
 sky130_fd_sc_hd__xnor2_4 _14161_ (.A(_06752_),
    .B(_06760_),
    .Y(net122));
 sky130_fd_sc_hd__and3_1 _14162_ (.A(_06730_),
    .B(_06731_),
    .C(_06732_),
    .X(_06761_));
 sky130_fd_sc_hd__and3_1 _14163_ (.A(_02742_),
    .B(_04013_),
    .C(_06702_),
    .X(_06762_));
 sky130_fd_sc_hd__xor2_1 _14164_ (.A(_06761_),
    .B(_06762_),
    .X(_06763_));
 sky130_fd_sc_hd__and2b_1 _14165_ (.A_N(_06708_),
    .B(_06735_),
    .X(_06764_));
 sky130_fd_sc_hd__or2_1 _14166_ (.A(_06764_),
    .B(_06741_),
    .X(_06766_));
 sky130_fd_sc_hd__xnor2_1 _14167_ (.A(_06763_),
    .B(_06766_),
    .Y(_06767_));
 sky130_fd_sc_hd__and3_1 _14168_ (.A(_06743_),
    .B(_06748_),
    .C(_06767_),
    .X(_06768_));
 sky130_fd_sc_hd__a21o_1 _14169_ (.A1(_06743_),
    .A2(_06748_),
    .B1(_06767_),
    .X(_06769_));
 sky130_fd_sc_hd__and2b_1 _14170_ (.A_N(_06768_),
    .B(_06769_),
    .X(_06770_));
 sky130_fd_sc_hd__xnor2_1 _14171_ (.A(_06750_),
    .B(_06770_),
    .Y(_06771_));
 sky130_fd_sc_hd__or4b_4 _14172_ (.A(_06616_),
    .B(_06642_),
    .C(_06753_),
    .D_N(_05841_),
    .X(_06772_));
 sky130_fd_sc_hd__or3b_1 _14173_ (.A(_06642_),
    .B(_06753_),
    .C_N(_06613_),
    .X(_06773_));
 sky130_fd_sc_hd__a2111o_1 _14174_ (.A1(_06772_),
    .A2(_06773_),
    .B1(_06636_),
    .C1(_06752_),
    .D1(_06759_),
    .X(_06774_));
 sky130_fd_sc_hd__xnor2_1 _14175_ (.A(_06771_),
    .B(_06774_),
    .Y(net123));
 sky130_fd_sc_hd__nor2_1 _14176_ (.A(_06752_),
    .B(_06759_),
    .Y(_06776_));
 sky130_fd_sc_hd__a21o_1 _14177_ (.A1(_05843_),
    .A2(_05849_),
    .B1(_06686_),
    .X(_06777_));
 sky130_fd_sc_hd__a21oi_4 _14178_ (.A1(_06687_),
    .A2(_06777_),
    .B1(_06645_),
    .Y(_06778_));
 sky130_fd_sc_hd__and2_1 _14179_ (.A(_06763_),
    .B(_06766_),
    .X(_06779_));
 sky130_fd_sc_hd__and4_1 _14180_ (.A(_02743_),
    .B(_04014_),
    .C(_02742_),
    .D(_04013_),
    .X(_06780_));
 sky130_fd_sc_hd__a211o_1 _14181_ (.A1(_06761_),
    .A2(_06762_),
    .B1(_06779_),
    .C1(_06780_),
    .X(_06781_));
 sky130_fd_sc_hd__inv_2 _14182_ (.A(_06770_),
    .Y(_06782_));
 sky130_fd_sc_hd__o21ai_1 _14183_ (.A1(_06750_),
    .A2(_06782_),
    .B1(_06769_),
    .Y(_06783_));
 sky130_fd_sc_hd__a311o_1 _14184_ (.A1(_06771_),
    .A2(_06776_),
    .A3(_06778_),
    .B1(_06781_),
    .C1(_06783_),
    .X(net124));
 sky130_fd_sc_hd__or4_1 _14185_ (.A(_05960_),
    .B(_06623_),
    .C(_06643_),
    .D(_06753_),
    .X(_06784_));
 sky130_fd_sc_hd__o32a_2 _14186_ (.A1(_06623_),
    .A2(_06643_),
    .A3(_06757_),
    .B1(_06784_),
    .B2(_05968_),
    .X(_06786_));
 sky130_fd_sc_hd__xnor2_4 _14187_ (.A(_06627_),
    .B(_06786_),
    .Y(net117));
 sky130_fd_sc_hd__nor2_2 _14188_ (.A(_06613_),
    .B(_06617_),
    .Y(_06787_));
 sky130_fd_sc_hd__xnor2_4 _14189_ (.A(_06787_),
    .B(_06620_),
    .Y(net110));
 sky130_fd_sc_hd__xor2_4 _14190_ (.A(_06632_),
    .B(_06689_),
    .X(net111));
 sky130_fd_sc_hd__xor2_4 _14191_ (.A(_06635_),
    .B(_06697_),
    .X(net112));
 sky130_fd_sc_hd__and3_1 _14192_ (.A(_06756_),
    .B(_06757_),
    .C(_06758_),
    .X(_06788_));
 sky130_fd_sc_hd__xnor2_1 _14193_ (.A(_06641_),
    .B(_06788_),
    .Y(net113));
 sky130_fd_sc_hd__and2_1 _14194_ (.A(_06772_),
    .B(_06773_),
    .X(_06789_));
 sky130_fd_sc_hd__xor2_1 _14195_ (.A(_06636_),
    .B(_06789_),
    .X(net114));
 sky130_fd_sc_hd__xnor2_4 _14196_ (.A(_06621_),
    .B(_06778_),
    .Y(net115));
 sky130_fd_sc_hd__or3_2 _14197_ (.A(_06621_),
    .B(_06644_),
    .C(_06697_),
    .X(_06791_));
 sky130_fd_sc_hd__xor2_4 _14198_ (.A(_06622_),
    .B(_06791_),
    .X(net116));
 sky130_fd_sc_hd__nor2_1 _14199_ (.A(_02357_),
    .B(_02390_),
    .Y(_06792_));
 sky130_fd_sc_hd__nor2_2 _14200_ (.A(_02401_),
    .B(_06792_),
    .Y(net120));
 sky130_fd_sc_hd__nand2_2 _14201_ (.A(_00344_),
    .B(_00410_),
    .Y(_06793_));
 sky130_fd_sc_hd__and2b_2 _14202_ (.A_N(_02938_),
    .B(_02927_),
    .X(_06794_));
 sky130_fd_sc_hd__xnor2_4 _14203_ (.A(_06793_),
    .B(_06794_),
    .Y(net127));
 sky130_fd_sc_hd__inv_2 _14204_ (.A(_02324_),
    .Y(_06795_));
 sky130_fd_sc_hd__nand2_2 _14205_ (.A(_02346_),
    .B(_06795_),
    .Y(_06796_));
 sky130_fd_sc_hd__xnor2_4 _14206_ (.A(_02270_),
    .B(_06796_),
    .Y(net109));
 sky130_fd_sc_hd__and2_1 _14207_ (.A(_01766_),
    .B(_01777_),
    .X(_06798_));
 sky130_fd_sc_hd__nor2_2 _14208_ (.A(_01788_),
    .B(_06798_),
    .Y(net98));
 sky130_fd_sc_hd__or2_1 _14209_ (.A(_01733_),
    .B(_01755_),
    .X(_06799_));
 sky130_fd_sc_hd__and2_1 _14210_ (.A(_01766_),
    .B(_06799_),
    .X(_06800_));
 sky130_fd_sc_hd__clkbuf_1 _14211_ (.A(_06800_),
    .X(net87));
 sky130_fd_sc_hd__a22oi_2 _14212_ (.A1(_00464_),
    .A2(_02138_),
    .B1(_00344_),
    .B2(_02051_),
    .Y(_06801_));
 sky130_fd_sc_hd__nor2_4 _14213_ (.A(_01755_),
    .B(_06801_),
    .Y(net76));
 sky130_fd_sc_hd__xor2_4 _14214_ (.A(net157),
    .B(_02423_),
    .X(net126));
 sky130_fd_sc_hd__xnor2_4 _14215_ (.A(_03642_),
    .B(_00229_),
    .Y(net66));
 sky130_fd_sc_hd__or2b_1 _14216_ (.A(_02412_),
    .B_N(_02248_),
    .X(_06803_));
 sky130_fd_sc_hd__xnor2_2 _14217_ (.A(_06803_),
    .B(_02401_),
    .Y(net125));
 sky130_fd_sc_hd__and2_1 _14218_ (.A(_00464_),
    .B(_00344_),
    .X(_06804_));
 sky130_fd_sc_hd__clkbuf_1 _14219_ (.A(_06804_),
    .X(net65));
 sky130_fd_sc_hd__inv_2 _14220_ (.A(_00404_),
    .Y(_06805_));
 sky130_fd_sc_hd__nand2_1 _14221_ (.A(_00405_),
    .B(_06805_),
    .Y(_06806_));
 sky130_fd_sc_hd__xnor2_2 _14222_ (.A(_00401_),
    .B(_06806_),
    .Y(net72));
 sky130_fd_sc_hd__and2_1 _14223_ (.A(_00406_),
    .B(_00408_),
    .X(_06807_));
 sky130_fd_sc_hd__nor2_1 _14224_ (.A(_00406_),
    .B(_00408_),
    .Y(_06808_));
 sky130_fd_sc_hd__nor2_2 _14225_ (.A(_06807_),
    .B(_06808_),
    .Y(net73));
 sky130_fd_sc_hd__xor2_2 _14226_ (.A(_00224_),
    .B(_00231_),
    .X(net67));
 sky130_fd_sc_hd__xor2_1 _14227_ (.A(_00233_),
    .B(_00241_),
    .X(net68));
 sky130_fd_sc_hd__mux2_4 _14228_ (.A0(_00244_),
    .A1(_00245_),
    .S(_00242_),
    .X(_06810_));
 sky130_fd_sc_hd__inv_2 _14229_ (.A(_06810_),
    .Y(net69));
 sky130_fd_sc_hd__xor2_4 _14230_ (.A(_00206_),
    .B(_00360_),
    .X(net70));
 sky130_fd_sc_hd__xnor2_1 _14231_ (.A(_00249_),
    .B(_00361_),
    .Y(net71));
 sky130_fd_sc_hd__or2b_1 _14232_ (.A(_00409_),
    .B_N(_00400_),
    .X(_06811_));
 sky130_fd_sc_hd__xnor2_2 _14233_ (.A(_06811_),
    .B(_06807_),
    .Y(net74));
 sky130_fd_sc_hd__buf_4 input1 (.A(a[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_4 input10 (.A(a[18]),
    .X(net10));
 sky130_fd_sc_hd__buf_4 input11 (.A(a[19]),
    .X(net11));
 sky130_fd_sc_hd__buf_12 input12 (.A(a[1]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_4 input13 (.A(a[20]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_4 input14 (.A(a[21]),
    .X(net14));
 sky130_fd_sc_hd__buf_4 input15 (.A(a[22]),
    .X(net15));
 sky130_fd_sc_hd__dlymetal6s2s_1 input16 (.A(a[23]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 input17 (.A(a[24]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(a[25]),
    .X(net18));
 sky130_fd_sc_hd__buf_4 input19 (.A(a[26]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(a[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_4 input20 (.A(a[27]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_4 input21 (.A(a[28]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_4 input22 (.A(a[29]),
    .X(net22));
 sky130_fd_sc_hd__buf_8 input23 (.A(a[2]),
    .X(net23));
 sky130_fd_sc_hd__buf_4 input24 (.A(a[30]),
    .X(net24));
 sky130_fd_sc_hd__buf_1 input25 (.A(a[31]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_4 input26 (.A(a[3]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_4 input27 (.A(a[4]),
    .X(net27));
 sky130_fd_sc_hd__buf_6 input28 (.A(a[5]),
    .X(net28));
 sky130_fd_sc_hd__buf_4 input29 (.A(a[6]),
    .X(net29));
 sky130_fd_sc_hd__buf_1 input3 (.A(a[11]),
    .X(net3));
 sky130_fd_sc_hd__buf_2 input30 (.A(a[7]),
    .X(net30));
 sky130_fd_sc_hd__buf_2 input31 (.A(a[8]),
    .X(net31));
 sky130_fd_sc_hd__buf_2 input32 (.A(a[9]),
    .X(net32));
 sky130_fd_sc_hd__buf_6 input33 (.A(b[0]),
    .X(net33));
 sky130_fd_sc_hd__buf_4 input34 (.A(b[10]),
    .X(net34));
 sky130_fd_sc_hd__buf_2 input35 (.A(b[11]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_4 input36 (.A(b[12]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_4 input37 (.A(b[13]),
    .X(net37));
 sky130_fd_sc_hd__buf_4 input38 (.A(b[14]),
    .X(net38));
 sky130_fd_sc_hd__buf_2 input39 (.A(b[15]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_8 input4 (.A(a[12]),
    .X(net4));
 sky130_fd_sc_hd__buf_4 input40 (.A(b[16]),
    .X(net40));
 sky130_fd_sc_hd__buf_1 input41 (.A(b[17]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_2 input42 (.A(b[18]),
    .X(net42));
 sky130_fd_sc_hd__buf_2 input43 (.A(b[19]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_8 input44 (.A(b[1]),
    .X(net44));
 sky130_fd_sc_hd__buf_4 input45 (.A(b[20]),
    .X(net45));
 sky130_fd_sc_hd__buf_4 input46 (.A(b[21]),
    .X(net46));
 sky130_fd_sc_hd__buf_4 input47 (.A(b[22]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_4 input48 (.A(b[23]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_4 input49 (.A(b[24]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_4 input5 (.A(a[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_4 input50 (.A(b[25]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_2 input51 (.A(b[26]),
    .X(net51));
 sky130_fd_sc_hd__buf_4 input52 (.A(b[27]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_2 input53 (.A(b[28]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_4 input54 (.A(b[29]),
    .X(net54));
 sky130_fd_sc_hd__buf_6 input55 (.A(b[2]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_4 input56 (.A(b[30]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_4 input57 (.A(b[31]),
    .X(net57));
 sky130_fd_sc_hd__buf_8 input58 (.A(b[3]),
    .X(net58));
 sky130_fd_sc_hd__buf_4 input59 (.A(b[4]),
    .X(net59));
 sky130_fd_sc_hd__buf_4 input6 (.A(a[14]),
    .X(net6));
 sky130_fd_sc_hd__buf_4 input60 (.A(b[5]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_4 input61 (.A(b[6]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_8 input62 (.A(b[7]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_8 input63 (.A(b[8]),
    .X(net63));
 sky130_fd_sc_hd__buf_4 input64 (.A(b[9]),
    .X(net64));
 sky130_fd_sc_hd__buf_4 input7 (.A(a[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_4 input8 (.A(a[16]),
    .X(net8));
 sky130_fd_sc_hd__buf_4 input9 (.A(a[17]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 max_cap1 (.A(_03504_),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_2 max_cap130 (.A(_05595_),
    .X(net130));
 sky130_fd_sc_hd__buf_1 max_cap132 (.A(_06562_),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_1 max_cap133 (.A(net134),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_1 max_cap134 (.A(_06504_),
    .X(net134));
 sky130_fd_sc_hd__buf_1 max_cap135 (.A(_06583_),
    .X(net135));
 sky130_fd_sc_hd__buf_1 max_cap138 (.A(_03504_),
    .X(net138));
 sky130_fd_sc_hd__buf_1 max_cap139 (.A(net180),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_2 max_cap140 (.A(_03455_),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_1 max_cap141 (.A(_06150_),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_1 max_cap142 (.A(_03701_),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_1 max_cap143 (.A(_01731_),
    .X(net143));
 sky130_fd_sc_hd__buf_1 max_cap144 (.A(_04299_),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_1 max_cap145 (.A(_00313_),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_1 max_cap146 (.A(_04265_),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_1 max_cap2 (.A(net180),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_4 output100 (.A(net100),
    .X(prod[41]));
 sky130_fd_sc_hd__clkbuf_4 output101 (.A(net101),
    .X(prod[42]));
 sky130_fd_sc_hd__clkbuf_4 output102 (.A(net102),
    .X(prod[43]));
 sky130_fd_sc_hd__clkbuf_4 output103 (.A(net103),
    .X(prod[44]));
 sky130_fd_sc_hd__clkbuf_4 output104 (.A(net104),
    .X(prod[45]));
 sky130_fd_sc_hd__clkbuf_4 output105 (.A(net105),
    .X(prod[46]));
 sky130_fd_sc_hd__clkbuf_4 output106 (.A(net106),
    .X(prod[47]));
 sky130_fd_sc_hd__clkbuf_4 output107 (.A(net107),
    .X(prod[48]));
 sky130_fd_sc_hd__clkbuf_4 output108 (.A(net108),
    .X(prod[49]));
 sky130_fd_sc_hd__clkbuf_4 output109 (.A(net109),
    .X(prod[4]));
 sky130_fd_sc_hd__clkbuf_4 output110 (.A(net110),
    .X(prod[50]));
 sky130_fd_sc_hd__clkbuf_4 output111 (.A(net111),
    .X(prod[51]));
 sky130_fd_sc_hd__clkbuf_4 output112 (.A(net112),
    .X(prod[52]));
 sky130_fd_sc_hd__clkbuf_4 output113 (.A(net129),
    .X(prod[53]));
 sky130_fd_sc_hd__clkbuf_4 output114 (.A(net114),
    .X(prod[54]));
 sky130_fd_sc_hd__buf_2 output115 (.A(net115),
    .X(prod[55]));
 sky130_fd_sc_hd__buf_4 output116 (.A(net116),
    .X(prod[56]));
 sky130_fd_sc_hd__clkbuf_4 output117 (.A(net117),
    .X(prod[57]));
 sky130_fd_sc_hd__clkbuf_4 output118 (.A(net118),
    .X(prod[58]));
 sky130_fd_sc_hd__buf_6 output119 (.A(net119),
    .X(prod[59]));
 sky130_fd_sc_hd__clkbuf_4 output120 (.A(net120),
    .X(prod[5]));
 sky130_fd_sc_hd__buf_6 output121 (.A(net121),
    .X(prod[60]));
 sky130_fd_sc_hd__buf_6 output122 (.A(net122),
    .X(prod[61]));
 sky130_fd_sc_hd__buf_4 output123 (.A(net123),
    .X(prod[62]));
 sky130_fd_sc_hd__clkbuf_4 output124 (.A(net124),
    .X(prod[63]));
 sky130_fd_sc_hd__clkbuf_4 output125 (.A(net125),
    .X(prod[6]));
 sky130_fd_sc_hd__clkbuf_4 output126 (.A(net126),
    .X(prod[7]));
 sky130_fd_sc_hd__clkbuf_4 output127 (.A(net127),
    .X(prod[8]));
 sky130_fd_sc_hd__buf_2 output128 (.A(net128),
    .X(prod[9]));
 sky130_fd_sc_hd__clkbuf_4 output65 (.A(net65),
    .X(prod[0]));
 sky130_fd_sc_hd__clkbuf_4 output66 (.A(net66),
    .X(prod[10]));
 sky130_fd_sc_hd__clkbuf_4 output67 (.A(net67),
    .X(prod[11]));
 sky130_fd_sc_hd__clkbuf_4 output68 (.A(net68),
    .X(prod[12]));
 sky130_fd_sc_hd__clkbuf_4 output69 (.A(net69),
    .X(prod[13]));
 sky130_fd_sc_hd__clkbuf_4 output70 (.A(net70),
    .X(prod[14]));
 sky130_fd_sc_hd__clkbuf_4 output71 (.A(net71),
    .X(prod[15]));
 sky130_fd_sc_hd__clkbuf_4 output72 (.A(net72),
    .X(prod[16]));
 sky130_fd_sc_hd__clkbuf_4 output73 (.A(net73),
    .X(prod[17]));
 sky130_fd_sc_hd__clkbuf_4 output74 (.A(net74),
    .X(prod[18]));
 sky130_fd_sc_hd__clkbuf_4 output75 (.A(net75),
    .X(prod[19]));
 sky130_fd_sc_hd__clkbuf_4 output76 (.A(net76),
    .X(prod[1]));
 sky130_fd_sc_hd__clkbuf_4 output77 (.A(net77),
    .X(prod[20]));
 sky130_fd_sc_hd__buf_2 output78 (.A(net78),
    .X(prod[21]));
 sky130_fd_sc_hd__clkbuf_4 output79 (.A(net79),
    .X(prod[22]));
 sky130_fd_sc_hd__clkbuf_4 output80 (.A(net80),
    .X(prod[23]));
 sky130_fd_sc_hd__clkbuf_4 output81 (.A(net81),
    .X(prod[24]));
 sky130_fd_sc_hd__clkbuf_4 output82 (.A(net82),
    .X(prod[25]));
 sky130_fd_sc_hd__clkbuf_4 output83 (.A(net83),
    .X(prod[26]));
 sky130_fd_sc_hd__clkbuf_4 output84 (.A(net84),
    .X(prod[27]));
 sky130_fd_sc_hd__clkbuf_4 output85 (.A(net85),
    .X(prod[28]));
 sky130_fd_sc_hd__clkbuf_4 output86 (.A(net86),
    .X(prod[29]));
 sky130_fd_sc_hd__buf_2 output87 (.A(net87),
    .X(prod[2]));
 sky130_fd_sc_hd__clkbuf_4 output88 (.A(net88),
    .X(prod[30]));
 sky130_fd_sc_hd__buf_2 output89 (.A(net89),
    .X(prod[31]));
 sky130_fd_sc_hd__clkbuf_4 output90 (.A(net90),
    .X(prod[32]));
 sky130_fd_sc_hd__clkbuf_4 output91 (.A(net91),
    .X(prod[33]));
 sky130_fd_sc_hd__clkbuf_4 output92 (.A(net92),
    .X(prod[34]));
 sky130_fd_sc_hd__clkbuf_4 output93 (.A(net93),
    .X(prod[35]));
 sky130_fd_sc_hd__buf_2 output94 (.A(net94),
    .X(prod[36]));
 sky130_fd_sc_hd__buf_2 output95 (.A(net95),
    .X(prod[37]));
 sky130_fd_sc_hd__clkbuf_4 output96 (.A(net96),
    .X(prod[38]));
 sky130_fd_sc_hd__buf_2 output97 (.A(net97),
    .X(prod[39]));
 sky130_fd_sc_hd__clkbuf_4 output98 (.A(net98),
    .X(prod[3]));
 sky130_fd_sc_hd__clkbuf_4 output99 (.A(net99),
    .X(prod[40]));
 sky130_fd_sc_hd__clkbuf_2 rebuffer1 (.A(_03235_),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_1 rebuffer10 (.A(_01799_),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_2 rebuffer11 (.A(_01985_),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_1 rebuffer12 (.A(_07060_),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_1 rebuffer13 (.A(_07060_),
    .X(net159));
 sky130_fd_sc_hd__buf_1 rebuffer14 (.A(_00588_),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_1 rebuffer15 (.A(_00716_),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_1 rebuffer16 (.A(net163),
    .X(net162));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer17 (.A(_00182_),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_1 rebuffer18 (.A(_04400_),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_2 rebuffer19 (.A(_07039_),
    .X(net165));
 sky130_fd_sc_hd__buf_1 rebuffer2 (.A(_06932_),
    .X(net148));
 sky130_fd_sc_hd__buf_1 rebuffer20 (.A(_06934_),
    .X(net166));
 sky130_fd_sc_hd__dlygate4sd3_1 rebuffer21 (.A(net183),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_1 rebuffer22 (.A(_01164_),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_1 rebuffer23 (.A(net168),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_1 rebuffer24 (.A(_04697_),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_1 rebuffer25 (.A(_07061_),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_1 rebuffer26 (.A(net171),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_1 rebuffer27 (.A(_07047_),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_1 rebuffer28 (.A(net173),
    .X(net174));
 sky130_fd_sc_hd__buf_1 rebuffer29 (.A(_00716_),
    .X(net175));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer3 (.A(_01810_),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_1 rebuffer30 (.A(_00923_),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_2 rebuffer31 (.A(_00923_),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_2 rebuffer32 (.A(_06065_),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_1 rebuffer33 (.A(_02083_),
    .X(net184));
 sky130_fd_sc_hd__dlymetal6s4s_1 rebuffer34 (.A(_04977_),
    .X(net185));
 sky130_fd_sc_hd__buf_6 rebuffer35 (.A(_04596_),
    .X(net186));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer36 (.A(_05967_),
    .X(net187));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer37 (.A(_03367_),
    .X(net188));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer38 (.A(_02740_),
    .X(net189));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer39 (.A(_05423_),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_1 rebuffer4 (.A(_06142_),
    .X(net150));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer40 (.A(_03246_),
    .X(net191));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer41 (.A(_03378_),
    .X(net192));
 sky130_fd_sc_hd__buf_1 rebuffer5 (.A(_05522_),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_2 rebuffer6 (.A(_02576_),
    .X(net152));
 sky130_fd_sc_hd__buf_1 rebuffer7 (.A(_00825_),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_1 rebuffer8 (.A(_04675_),
    .X(net154));
 sky130_fd_sc_hd__buf_1 rebuffer9 (.A(_05037_),
    .X(net155));
 sky130_fd_sc_hd__buf_6 split17 (.A(_00716_),
    .X(net163));
 sky130_fd_sc_hd__buf_2 split3 (.A(_00869_),
    .X(net149));
 sky130_fd_sc_hd__buf_4 wire129 (.A(net113),
    .X(net129));
 sky130_fd_sc_hd__buf_2 wire131 (.A(_01242_),
    .X(net131));
 sky130_fd_sc_hd__buf_1 wire136 (.A(_06487_),
    .X(net136));
 sky130_fd_sc_hd__buf_1 wire137 (.A(_06364_),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_1 wire3 (.A(_06691_),
    .X(net180));
endmodule

